`timescale 1ns / 1ps

module gif (input clock, input [6:0] x, y, input [2:0] machine_state, output reg [15:0] oled_data = 0);
	reg [4:0]frame_rate = 5'd3;
	reg [3:0]frame_no = 4'd1;
	reg [31:0]COUNT = 32'b1;
	reg slow_clk = 1'b0;

	always @ (*) begin
		if (machine_state == 3'd6) begin
			case ({frame_no, x, y})
				18'b000100011000001000: oled_data = 16'b1001110000001011;
				18'b000100011010001000: oled_data = 16'b1010010000101100;
				18'b000100011100001000: oled_data = 16'b1010010000101100;
				18'b000100011110001000: oled_data = 16'b1010110000101011;
				18'b000100100000001000: oled_data = 16'b1010110000101011;
				18'b000100100010001000: oled_data = 16'b1010110000101011;
				18'b000100100100001000: oled_data = 16'b1010110000101011;
				18'b000100100110001000: oled_data = 16'b1010110000101011;
				18'b000100101000001000: oled_data = 16'b1010010000001011;
				18'b000100101010001000: oled_data = 16'b1101111000010111;
				18'b000100101100001000: oled_data = 16'b1110110111011000;
				18'b000100101110001000: oled_data = 16'b1110010011010110;
				18'b000100110000001000: oled_data = 16'b1110010011010110;
				18'b000100110010001000: oled_data = 16'b1110010010110110;
				18'b000100110100001000: oled_data = 16'b1110010010110110;
				18'b000100110110001000: oled_data = 16'b1110010010110110;
				18'b000100111000001000: oled_data = 16'b1110010010110110;
				18'b000100111010001000: oled_data = 16'b1110010010110110;
				18'b000100111100001000: oled_data = 16'b1110010010110110;
				18'b000100111110001000: oled_data = 16'b1110010010110110;
				18'b000101000000001000: oled_data = 16'b1110010010110110;
				18'b000101000010001000: oled_data = 16'b1110010010110110;
				18'b000101000100001000: oled_data = 16'b1110010010110110;
				18'b000101000110001000: oled_data = 16'b1110010010110110;
				18'b000101001000001000: oled_data = 16'b1110010010110110;
				18'b000101001010001000: oled_data = 16'b1110010010110110;
				18'b000101001100001000: oled_data = 16'b1110010010110110;
				18'b000101001110001000: oled_data = 16'b1110010010110110;
				18'b000101010000001000: oled_data = 16'b1110010010110110;
				18'b000101010010001000: oled_data = 16'b1110010010110110;
				18'b000101010100001000: oled_data = 16'b1110010010110110;
				18'b000101010110001000: oled_data = 16'b1110010010110110;
				18'b000101011000001000: oled_data = 16'b1110010010110110;
				18'b000101011010001000: oled_data = 16'b1110010011010110;
				18'b000101011100001000: oled_data = 16'b1101110010110101;
				18'b000101011110001000: oled_data = 16'b1110010010110110;
				18'b000101100000001000: oled_data = 16'b1110010011010110;
				18'b000101100010001000: oled_data = 16'b1110010010110110;
				18'b000101100100001000: oled_data = 16'b1110010010110110;
				18'b000101100110001000: oled_data = 16'b1101110011010101;
				18'b000101101000001000: oled_data = 16'b1101010010010100;
				18'b000101101010001000: oled_data = 16'b1101110010010101;
				18'b000101101100001000: oled_data = 16'b1110010011110110;
				18'b000101101110001000: oled_data = 16'b1110010011010110;
				18'b000101110000001000: oled_data = 16'b1101110011010110;
				18'b000101110010001000: oled_data = 16'b1110010011110110;
				18'b000101110100001000: oled_data = 16'b1101110011010110;
				18'b000101110110001000: oled_data = 16'b1101110011010101;
				18'b000101111000001000: oled_data = 16'b1101110011010101;
				18'b000101111010001000: oled_data = 16'b1101110010110101;
				18'b000101111100001000: oled_data = 16'b1101010001110100;
				18'b000101111110001000: oled_data = 16'b1101110011010101;
				18'b000110000000001000: oled_data = 16'b1101110011010110;
				18'b000110000010001000: oled_data = 16'b1101110011010110;
				18'b000110000100001000: oled_data = 16'b1101010011110101;
				18'b000110000110001000: oled_data = 16'b1110111001111011;
				18'b000110001000001000: oled_data = 16'b1110011000111001;
				18'b000110001010001000: oled_data = 16'b0111001010101000;
				18'b000110001100001000: oled_data = 16'b0110101010100101;
				18'b000110001110001000: oled_data = 16'b0111101100000111;
				18'b000110010000001000: oled_data = 16'b0111101100000111;
				18'b000110010010001000: oled_data = 16'b0111101011100111;
				18'b000110010100001000: oled_data = 16'b0111101100000111;
				18'b000110010110001000: oled_data = 16'b0111001011101000;
				18'b000110011000001000: oled_data = 16'b0110101011001000;
				18'b000110011010001000: oled_data = 16'b0110101011001000;
				18'b000110011100001000: oled_data = 16'b0110001010101000;
				18'b000110011110001000: oled_data = 16'b0101101010000111;
				18'b000110100000001000: oled_data = 16'b0101101010001000;
				18'b000110100010001000: oled_data = 16'b0101001001101000;
				18'b000110100100001000: oled_data = 16'b0101001001101000;
				18'b000110100110001000: oled_data = 16'b0101001001101000;
				18'b000100011000001001: oled_data = 16'b1011010001101011;
				18'b000100011010001001: oled_data = 16'b1011010001001011;
				18'b000100011100001001: oled_data = 16'b1011010001001011;
				18'b000100011110001001: oled_data = 16'b1011010001001011;
				18'b000100100000001001: oled_data = 16'b1011010001001011;
				18'b000100100010001001: oled_data = 16'b1011010001001011;
				18'b000100100100001001: oled_data = 16'b1011010001001011;
				18'b000100100110001001: oled_data = 16'b1010110000101010;
				18'b000100101000001001: oled_data = 16'b1100010100010001;
				18'b000100101010001001: oled_data = 16'b1111011001011010;
				18'b000100101100001001: oled_data = 16'b1101110011110110;
				18'b000100101110001001: oled_data = 16'b1101110011010101;
				18'b000100110000001001: oled_data = 16'b1101010010010100;
				18'b000100110010001001: oled_data = 16'b1101110011010101;
				18'b000100110100001001: oled_data = 16'b1101110011010101;
				18'b000100110110001001: oled_data = 16'b1101110011010101;
				18'b000100111000001001: oled_data = 16'b1101110011010101;
				18'b000100111010001001: oled_data = 16'b1101110011010101;
				18'b000100111100001001: oled_data = 16'b1101110011010101;
				18'b000100111110001001: oled_data = 16'b1101110011010101;
				18'b000101000000001001: oled_data = 16'b1101110011010101;
				18'b000101000010001001: oled_data = 16'b1101110011010101;
				18'b000101000100001001: oled_data = 16'b1101110011010101;
				18'b000101000110001001: oled_data = 16'b1101110011010101;
				18'b000101001000001001: oled_data = 16'b1101110011010101;
				18'b000101001010001001: oled_data = 16'b1101110011010101;
				18'b000101001100001001: oled_data = 16'b1101110011010101;
				18'b000101001110001001: oled_data = 16'b1101110011010101;
				18'b000101010000001001: oled_data = 16'b1101110011010101;
				18'b000101010010001001: oled_data = 16'b1101110011010101;
				18'b000101010100001001: oled_data = 16'b1101110011010101;
				18'b000101010110001001: oled_data = 16'b1101110011010101;
				18'b000101011000001001: oled_data = 16'b1101110011010101;
				18'b000101011010001001: oled_data = 16'b1101110011010101;
				18'b000101011100001001: oled_data = 16'b1101110010010101;
				18'b000101011110001001: oled_data = 16'b1101010001110100;
				18'b000101100000001001: oled_data = 16'b1101110010110101;
				18'b000101100010001001: oled_data = 16'b1101110011010101;
				18'b000101100100001001: oled_data = 16'b1101110011010101;
				18'b000101100110001001: oled_data = 16'b1101110011010101;
				18'b000101101000001001: oled_data = 16'b1101110011010110;
				18'b000101101010001001: oled_data = 16'b1101010001110100;
				18'b000101101100001001: oled_data = 16'b1101010010010101;
				18'b000101101110001001: oled_data = 16'b1101110011010110;
				18'b000101110000001001: oled_data = 16'b1101110011010101;
				18'b000101110010001001: oled_data = 16'b1101110011010110;
				18'b000101110100001001: oled_data = 16'b1110010011110110;
				18'b000101110110001001: oled_data = 16'b1101110011010101;
				18'b000101111000001001: oled_data = 16'b1101110011010101;
				18'b000101111010001001: oled_data = 16'b1101110011010110;
				18'b000101111100001001: oled_data = 16'b1101010010010100;
				18'b000101111110001001: oled_data = 16'b1101010010010100;
				18'b000110000000001001: oled_data = 16'b1101110011010101;
				18'b000110000010001001: oled_data = 16'b1101110011010101;
				18'b000110000100001001: oled_data = 16'b1101110011110101;
				18'b000110000110001001: oled_data = 16'b1101010100110110;
				18'b000110001000001001: oled_data = 16'b1111011011011100;
				18'b000110001010001001: oled_data = 16'b1001110000101110;
				18'b000110001100001001: oled_data = 16'b0111001011000110;
				18'b000110001110001001: oled_data = 16'b0111001011000111;
				18'b000110010000001001: oled_data = 16'b1000001100101000;
				18'b000110010010001001: oled_data = 16'b1000001100101000;
				18'b000110010100001001: oled_data = 16'b1000001100101000;
				18'b000110010110001001: oled_data = 16'b1000001101001000;
				18'b000110011000001001: oled_data = 16'b1000101101001000;
				18'b000110011010001001: oled_data = 16'b1000101101101000;
				18'b000110011100001001: oled_data = 16'b1000101110001001;
				18'b000110011110001001: oled_data = 16'b1000101110001000;
				18'b000110100000001001: oled_data = 16'b1000101110101001;
				18'b000110100010001001: oled_data = 16'b0101101010101000;
				18'b000110100100001001: oled_data = 16'b0100001000001000;
				18'b000110100110001001: oled_data = 16'b0100001000101000;
				18'b000100011000001010: oled_data = 16'b1011010001101011;
				18'b000100011010001010: oled_data = 16'b1011010001101011;
				18'b000100011100001010: oled_data = 16'b1010110001001011;
				18'b000100011110001010: oled_data = 16'b1010110001001011;
				18'b000100100000001010: oled_data = 16'b1010010000101011;
				18'b000100100010001010: oled_data = 16'b1001101111101010;
				18'b000100100100001010: oled_data = 16'b1001001110101001;
				18'b000100100110001010: oled_data = 16'b1001001110101010;
				18'b000100101000001010: oled_data = 16'b1110011000111000;
				18'b000100101010001010: oled_data = 16'b1110010101010111;
				18'b000100101100001010: oled_data = 16'b1110010011010101;
				18'b000100101110001010: oled_data = 16'b1101010001110100;
				18'b000100110000001010: oled_data = 16'b1101110010110101;
				18'b000100110010001010: oled_data = 16'b1101110011010101;
				18'b000100110100001010: oled_data = 16'b1101110011010101;
				18'b000100110110001010: oled_data = 16'b1101110011010101;
				18'b000100111000001010: oled_data = 16'b1101110011010101;
				18'b000100111010001010: oled_data = 16'b1101110011010101;
				18'b000100111100001010: oled_data = 16'b1101110011010101;
				18'b000100111110001010: oled_data = 16'b1101110011010101;
				18'b000101000000001010: oled_data = 16'b1101110011010101;
				18'b000101000010001010: oled_data = 16'b1101110011010101;
				18'b000101000100001010: oled_data = 16'b1101110011010101;
				18'b000101000110001010: oled_data = 16'b1101110011010101;
				18'b000101001000001010: oled_data = 16'b1101110011010101;
				18'b000101001010001010: oled_data = 16'b1101110011010101;
				18'b000101001100001010: oled_data = 16'b1101110011010101;
				18'b000101001110001010: oled_data = 16'b1101110011010101;
				18'b000101010000001010: oled_data = 16'b1101110011010101;
				18'b000101010010001010: oled_data = 16'b1101110011010101;
				18'b000101010100001010: oled_data = 16'b1101110011010101;
				18'b000101010110001010: oled_data = 16'b1101110011010101;
				18'b000101011000001010: oled_data = 16'b1101110011010101;
				18'b000101011010001010: oled_data = 16'b1101110011010101;
				18'b000101011100001010: oled_data = 16'b1101110011010101;
				18'b000101011110001010: oled_data = 16'b1101110010110101;
				18'b000101100000001010: oled_data = 16'b1101010001110100;
				18'b000101100010001010: oled_data = 16'b1101110010110101;
				18'b000101100100001010: oled_data = 16'b1101110011010101;
				18'b000101100110001010: oled_data = 16'b1101110011010101;
				18'b000101101000001010: oled_data = 16'b1101110011010110;
				18'b000101101010001010: oled_data = 16'b1101110011010101;
				18'b000101101100001010: oled_data = 16'b1101010010010100;
				18'b000101101110001010: oled_data = 16'b1101010001110100;
				18'b000101110000001010: oled_data = 16'b1101110011010110;
				18'b000101110010001010: oled_data = 16'b1101110011010101;
				18'b000101110100001010: oled_data = 16'b1110010011010110;
				18'b000101110110001010: oled_data = 16'b1110010011010110;
				18'b000101111000001010: oled_data = 16'b1101110011010101;
				18'b000101111010001010: oled_data = 16'b1101110011010101;
				18'b000101111100001010: oled_data = 16'b1101110011010110;
				18'b000101111110001010: oled_data = 16'b1101010001110100;
				18'b000110000000001010: oled_data = 16'b1101110011010101;
				18'b000110000010001010: oled_data = 16'b1101110011010101;
				18'b000110000100001010: oled_data = 16'b1101110011110110;
				18'b000110000110001010: oled_data = 16'b1101010011010101;
				18'b000110001000001010: oled_data = 16'b1110011000111001;
				18'b000110001010001010: oled_data = 16'b1100110110110110;
				18'b000110001100001010: oled_data = 16'b0100000111100110;
				18'b000110001110001010: oled_data = 16'b0101001000000110;
				18'b000110010000001010: oled_data = 16'b0110001001100111;
				18'b000110010010001010: oled_data = 16'b0111001010100111;
				18'b000110010100001010: oled_data = 16'b0111101011101000;
				18'b000110010110001010: oled_data = 16'b1000001100101000;
				18'b000110011000001010: oled_data = 16'b1000001101001000;
				18'b000110011010001010: oled_data = 16'b1000101101101000;
				18'b000110011100001010: oled_data = 16'b1001001101101000;
				18'b000110011110001010: oled_data = 16'b1000101101101000;
				18'b000110100000001010: oled_data = 16'b1000101101101001;
				18'b000110100010001010: oled_data = 16'b0111101011101010;
				18'b000110100100001010: oled_data = 16'b1001001101001101;
				18'b000110100110001010: oled_data = 16'b1011010000010000;
				18'b000100011000001011: oled_data = 16'b1001001111101010;
				18'b000100011010001011: oled_data = 16'b1000101110001001;
				18'b000100011100001011: oled_data = 16'b0111101100101001;
				18'b000100011110001011: oled_data = 16'b0110101011101001;
				18'b000100100000001011: oled_data = 16'b0110001010101001;
				18'b000100100010001011: oled_data = 16'b0101101001101000;
				18'b000100100100001011: oled_data = 16'b0101101001001000;
				18'b000100100110001011: oled_data = 16'b1001110001010000;
				18'b000100101000001011: oled_data = 16'b1110111001011010;
				18'b000100101010001011: oled_data = 16'b1101110011010101;
				18'b000100101100001011: oled_data = 16'b1101110010110101;
				18'b000100101110001011: oled_data = 16'b1101010010010100;
				18'b000100110000001011: oled_data = 16'b1110010011110110;
				18'b000100110010001011: oled_data = 16'b1101110011010110;
				18'b000100110100001011: oled_data = 16'b1101110011010101;
				18'b000100110110001011: oled_data = 16'b1101110011010110;
				18'b000100111000001011: oled_data = 16'b1101110011010110;
				18'b000100111010001011: oled_data = 16'b1101110011010110;
				18'b000100111100001011: oled_data = 16'b1101110011010110;
				18'b000100111110001011: oled_data = 16'b1101110011010110;
				18'b000101000000001011: oled_data = 16'b1101110011010110;
				18'b000101000010001011: oled_data = 16'b1101110011010110;
				18'b000101000100001011: oled_data = 16'b1101110011010110;
				18'b000101000110001011: oled_data = 16'b1101110011010110;
				18'b000101001000001011: oled_data = 16'b1101110011010110;
				18'b000101001010001011: oled_data = 16'b1101110011010110;
				18'b000101001100001011: oled_data = 16'b1101110011010110;
				18'b000101001110001011: oled_data = 16'b1101110011010110;
				18'b000101010000001011: oled_data = 16'b1101110011010110;
				18'b000101010010001011: oled_data = 16'b1101110011010110;
				18'b000101010100001011: oled_data = 16'b1101110011010110;
				18'b000101010110001011: oled_data = 16'b1101110011010110;
				18'b000101011000001011: oled_data = 16'b1101110011010110;
				18'b000101011010001011: oled_data = 16'b1101110011010110;
				18'b000101011100001011: oled_data = 16'b1101110011010110;
				18'b000101011110001011: oled_data = 16'b1101110011010110;
				18'b000101100000001011: oled_data = 16'b1101110010110101;
				18'b000101100010001011: oled_data = 16'b1101010001110100;
				18'b000101100100001011: oled_data = 16'b1101110010110101;
				18'b000101100110001011: oled_data = 16'b1101110011010101;
				18'b000101101000001011: oled_data = 16'b1110010101010111;
				18'b000101101010001011: oled_data = 16'b1110010100110111;
				18'b000101101100001011: oled_data = 16'b1110010011010110;
				18'b000101101110001011: oled_data = 16'b1100110001010011;
				18'b000101110000001011: oled_data = 16'b1100110000110011;
				18'b000101110010001011: oled_data = 16'b1110010011010110;
				18'b000101110100001011: oled_data = 16'b1101110011010110;
				18'b000101110110001011: oled_data = 16'b1101110011010101;
				18'b000101111000001011: oled_data = 16'b1101110011010101;
				18'b000101111010001011: oled_data = 16'b1101110011010110;
				18'b000101111100001011: oled_data = 16'b1101110011010110;
				18'b000101111110001011: oled_data = 16'b1101110010110101;
				18'b000110000000001011: oled_data = 16'b1101010001110100;
				18'b000110000010001011: oled_data = 16'b1101110011010110;
				18'b000110000100001011: oled_data = 16'b1101110011010110;
				18'b000110000110001011: oled_data = 16'b1101010010110101;
				18'b000110001000001011: oled_data = 16'b1101010011110101;
				18'b000110001010001011: oled_data = 16'b1110011001111010;
				18'b000110001100001011: oled_data = 16'b0101001001001001;
				18'b000110001110001011: oled_data = 16'b0010000101000101;
				18'b000110010000001011: oled_data = 16'b0010100101100110;
				18'b000110010010001011: oled_data = 16'b0010100110000110;
				18'b000110010100001011: oled_data = 16'b0011100111000111;
				18'b000110010110001011: oled_data = 16'b0100000111100111;
				18'b000110011000001011: oled_data = 16'b0100101000100111;
				18'b000110011010001011: oled_data = 16'b0101101001100110;
				18'b000110011100001011: oled_data = 16'b0111001011001000;
				18'b000110011110001011: oled_data = 16'b1010001110001011;
				18'b000110100000001011: oled_data = 16'b1100010001010000;
				18'b000110100010001011: oled_data = 16'b1101110010110010;
				18'b000110100100001011: oled_data = 16'b1110010001010001;
				18'b000110100110001011: oled_data = 16'b1100101101101110;
				18'b000100011000001100: oled_data = 16'b0101101010101000;
				18'b000100011010001100: oled_data = 16'b0110001010101000;
				18'b000100011100001100: oled_data = 16'b0110101011101010;
				18'b000100011110001100: oled_data = 16'b0111001100101010;
				18'b000100100000001100: oled_data = 16'b1000001101001010;
				18'b000100100010001100: oled_data = 16'b1000101110101011;
				18'b000100100100001100: oled_data = 16'b1001001111001011;
				18'b000100100110001100: oled_data = 16'b1101110111110111;
				18'b000100101000001100: oled_data = 16'b1101110101010111;
				18'b000100101010001100: oled_data = 16'b1101110011010110;
				18'b000100101100001100: oled_data = 16'b1101010010010100;
				18'b000100101110001100: oled_data = 16'b1101110011010101;
				18'b000100110000001100: oled_data = 16'b1110010011010110;
				18'b000100110010001100: oled_data = 16'b1101110011010110;
				18'b000100110100001100: oled_data = 16'b1101110011010101;
				18'b000100110110001100: oled_data = 16'b1101110011010110;
				18'b000100111000001100: oled_data = 16'b1101110011010110;
				18'b000100111010001100: oled_data = 16'b1101110011010110;
				18'b000100111100001100: oled_data = 16'b1101110011010110;
				18'b000100111110001100: oled_data = 16'b1101110011010110;
				18'b000101000000001100: oled_data = 16'b1101110011010110;
				18'b000101000010001100: oled_data = 16'b1101110011010110;
				18'b000101000100001100: oled_data = 16'b1101110011010110;
				18'b000101000110001100: oled_data = 16'b1101110011010110;
				18'b000101001000001100: oled_data = 16'b1101110011010110;
				18'b000101001010001100: oled_data = 16'b1101110010010101;
				18'b000101001100001100: oled_data = 16'b1101110010110101;
				18'b000101001110001100: oled_data = 16'b1101110011010110;
				18'b000101010000001100: oled_data = 16'b1101110011010110;
				18'b000101010010001100: oled_data = 16'b1101110011010110;
				18'b000101010100001100: oled_data = 16'b1101110011010110;
				18'b000101010110001100: oled_data = 16'b1101110011010110;
				18'b000101011000001100: oled_data = 16'b1101110011010110;
				18'b000101011010001100: oled_data = 16'b1101110011010110;
				18'b000101011100001100: oled_data = 16'b1101110011010110;
				18'b000101011110001100: oled_data = 16'b1101110011010110;
				18'b000101100000001100: oled_data = 16'b1101110011010101;
				18'b000101100010001100: oled_data = 16'b1101110010110101;
				18'b000101100100001100: oled_data = 16'b1100010000110011;
				18'b000101100110001100: oled_data = 16'b1101010010110101;
				18'b000101101000001100: oled_data = 16'b1101110100010110;
				18'b000101101010001100: oled_data = 16'b1110010101010111;
				18'b000101101100001100: oled_data = 16'b1110010011010110;
				18'b000101101110001100: oled_data = 16'b1110010011110110;
				18'b000101110000001100: oled_data = 16'b1100001111110010;
				18'b000101110010001100: oled_data = 16'b1100010000010010;
				18'b000101110100001100: oled_data = 16'b1110010011010110;
				18'b000101110110001100: oled_data = 16'b1101110011010101;
				18'b000101111000001100: oled_data = 16'b1101110011010101;
				18'b000101111010001100: oled_data = 16'b1101110011010110;
				18'b000101111100001100: oled_data = 16'b1101110011010101;
				18'b000101111110001100: oled_data = 16'b1101110011010110;
				18'b000110000000001100: oled_data = 16'b1101010001010100;
				18'b000110000010001100: oled_data = 16'b1101110011010101;
				18'b000110000100001100: oled_data = 16'b1101110011010110;
				18'b000110000110001100: oled_data = 16'b1101110010110101;
				18'b000110001000001100: oled_data = 16'b1101010010010100;
				18'b000110001010001100: oled_data = 16'b1110110110111000;
				18'b000110001100001100: oled_data = 16'b1000101111010000;
				18'b000110001110001100: oled_data = 16'b0010000100100101;
				18'b000110010000001100: oled_data = 16'b0010000101100110;
				18'b000110010010001100: oled_data = 16'b0010000101100110;
				18'b000110010100001100: oled_data = 16'b0010100110000111;
				18'b000110010110001100: oled_data = 16'b0010100110000111;
				18'b000110011000001100: oled_data = 16'b0011000110000110;
				18'b000110011010001100: oled_data = 16'b0111001010101010;
				18'b000110011100001100: oled_data = 16'b1011110001010001;
				18'b000110011110001100: oled_data = 16'b1110010011110100;
				18'b000110100000001100: oled_data = 16'b1101110000110001;
				18'b000110100010001100: oled_data = 16'b1100001100001101;
				18'b000110100100001100: oled_data = 16'b1010101001001001;
				18'b000110100110001100: oled_data = 16'b1010101000001000;
				18'b000100011000001101: oled_data = 16'b1001110000001011;
				18'b000100011010001101: oled_data = 16'b1010010000101010;
				18'b000100011100001101: oled_data = 16'b1010110000101011;
				18'b000100011110001101: oled_data = 16'b1010110000101011;
				18'b000100100000001101: oled_data = 16'b1010110000101011;
				18'b000100100010001101: oled_data = 16'b1010110000001011;
				18'b000100100100001101: oled_data = 16'b1011010010001110;
				18'b000100100110001101: oled_data = 16'b1110011000011000;
				18'b000100101000001101: oled_data = 16'b1101110011010110;
				18'b000100101010001101: oled_data = 16'b1101110011010101;
				18'b000100101100001101: oled_data = 16'b1101010001110100;
				18'b000100101110001101: oled_data = 16'b1110010011010110;
				18'b000100110000001101: oled_data = 16'b1101110011010110;
				18'b000100110010001101: oled_data = 16'b1101110011010110;
				18'b000100110100001101: oled_data = 16'b1101110011010110;
				18'b000100110110001101: oled_data = 16'b1101110010110101;
				18'b000100111000001101: oled_data = 16'b1101110010110101;
				18'b000100111010001101: oled_data = 16'b1101110011010101;
				18'b000100111100001101: oled_data = 16'b1101110011010101;
				18'b000100111110001101: oled_data = 16'b1101110011010101;
				18'b000101000000001101: oled_data = 16'b1101110011010101;
				18'b000101000010001101: oled_data = 16'b1101110011010101;
				18'b000101000100001101: oled_data = 16'b1101110011010101;
				18'b000101000110001101: oled_data = 16'b1101110011010101;
				18'b000101001000001101: oled_data = 16'b1101110011010110;
				18'b000101001010001101: oled_data = 16'b1101010010010100;
				18'b000101001100001101: oled_data = 16'b1101110010110101;
				18'b000101001110001101: oled_data = 16'b1101110011010101;
				18'b000101010000001101: oled_data = 16'b1101110011010101;
				18'b000101010010001101: oled_data = 16'b1101110011010101;
				18'b000101010100001101: oled_data = 16'b1101110011010101;
				18'b000101010110001101: oled_data = 16'b1101110011010101;
				18'b000101011000001101: oled_data = 16'b1101110011010101;
				18'b000101011010001101: oled_data = 16'b1101110011010101;
				18'b000101011100001101: oled_data = 16'b1101110011010101;
				18'b000101011110001101: oled_data = 16'b1101110011010101;
				18'b000101100000001101: oled_data = 16'b1101110011010101;
				18'b000101100010001101: oled_data = 16'b1101110011010110;
				18'b000101100100001101: oled_data = 16'b1101010010010100;
				18'b000101100110001101: oled_data = 16'b1100010000110011;
				18'b000101101000001101: oled_data = 16'b1101110011010101;
				18'b000101101010001101: oled_data = 16'b1101110011110110;
				18'b000101101100001101: oled_data = 16'b1110010011010110;
				18'b000101101110001101: oled_data = 16'b1110010011010110;
				18'b000101110000001101: oled_data = 16'b1101110011010101;
				18'b000101110010001101: oled_data = 16'b1011101110010001;
				18'b000101110100001101: oled_data = 16'b1100110000010011;
				18'b000101110110001101: oled_data = 16'b1110010011010110;
				18'b000101111000001101: oled_data = 16'b1101110011010101;
				18'b000101111010001101: oled_data = 16'b1101110011010101;
				18'b000101111100001101: oled_data = 16'b1101110011010101;
				18'b000101111110001101: oled_data = 16'b1101110011010110;
				18'b000110000000001101: oled_data = 16'b1101110010010101;
				18'b000110000010001101: oled_data = 16'b1101010010010100;
				18'b000110000100001101: oled_data = 16'b1101110011010110;
				18'b000110000110001101: oled_data = 16'b1101110011010101;
				18'b000110001000001101: oled_data = 16'b1101010001110100;
				18'b000110001010001101: oled_data = 16'b1101110011110110;
				18'b000110001100001101: oled_data = 16'b1010110011110100;
				18'b000110001110001101: oled_data = 16'b0010000100100101;
				18'b000110010000001101: oled_data = 16'b0010000101000110;
				18'b000110010010001101: oled_data = 16'b0010000101100110;
				18'b000110010100001101: oled_data = 16'b0010000101100110;
				18'b000110010110001101: oled_data = 16'b0100000111101000;
				18'b000110011000001101: oled_data = 16'b1010001111110000;
				18'b000110011010001101: oled_data = 16'b1110010011110100;
				18'b000110011100001101: oled_data = 16'b1101110010010010;
				18'b000110011110001101: oled_data = 16'b1100101101001101;
				18'b000110100000001101: oled_data = 16'b1011001001001001;
				18'b000110100010001101: oled_data = 16'b1011001000101001;
				18'b000110100100001101: oled_data = 16'b1010101000101000;
				18'b000110100110001101: oled_data = 16'b1010101000101000;
				18'b000100011000001110: oled_data = 16'b1010110001001011;
				18'b000100011010001110: oled_data = 16'b1010110001001011;
				18'b000100011100001110: oled_data = 16'b1011010001001011;
				18'b000100011110001110: oled_data = 16'b1010110000101011;
				18'b000100100000001110: oled_data = 16'b1010110000101011;
				18'b000100100010001110: oled_data = 16'b1010110000001011;
				18'b000100100100001110: oled_data = 16'b1100010100110010;
				18'b000100100110001110: oled_data = 16'b1110010110010111;
				18'b000100101000001110: oled_data = 16'b1101110011010110;
				18'b000100101010001110: oled_data = 16'b1101010010010101;
				18'b000100101100001110: oled_data = 16'b1101110010110101;
				18'b000100101110001110: oled_data = 16'b1101110011010101;
				18'b000100110000001110: oled_data = 16'b1101110011010110;
				18'b000100110010001110: oled_data = 16'b1101110011010110;
				18'b000100110100001110: oled_data = 16'b1101110011010101;
				18'b000100110110001110: oled_data = 16'b1101010001110100;
				18'b000100111000001110: oled_data = 16'b1101110011010101;
				18'b000100111010001110: oled_data = 16'b1101110011010110;
				18'b000100111100001110: oled_data = 16'b1101110011010101;
				18'b000100111110001110: oled_data = 16'b1101110011010101;
				18'b000101000000001110: oled_data = 16'b1101110011010101;
				18'b000101000010001110: oled_data = 16'b1101110010110101;
				18'b000101000100001110: oled_data = 16'b1101010010010100;
				18'b000101000110001110: oled_data = 16'b1101110011010110;
				18'b000101001000001110: oled_data = 16'b1101110011010110;
				18'b000101001010001110: oled_data = 16'b1101110010110101;
				18'b000101001100001110: oled_data = 16'b1101010010010101;
				18'b000101001110001110: oled_data = 16'b1101110011010110;
				18'b000101010000001110: oled_data = 16'b1101110011010101;
				18'b000101010010001110: oled_data = 16'b1101110011010101;
				18'b000101010100001110: oled_data = 16'b1101110011010101;
				18'b000101010110001110: oled_data = 16'b1101110011010101;
				18'b000101011000001110: oled_data = 16'b1101110011010101;
				18'b000101011010001110: oled_data = 16'b1101110011010101;
				18'b000101011100001110: oled_data = 16'b1101110011010101;
				18'b000101011110001110: oled_data = 16'b1101110011010101;
				18'b000101100000001110: oled_data = 16'b1101110011010101;
				18'b000101100010001110: oled_data = 16'b1101110011010101;
				18'b000101100100001110: oled_data = 16'b1101110011010110;
				18'b000101100110001110: oled_data = 16'b1101010010010100;
				18'b000101101000001110: oled_data = 16'b1100110001110011;
				18'b000101101010001110: oled_data = 16'b1101110010110101;
				18'b000101101100001110: oled_data = 16'b1110010011010110;
				18'b000101101110001110: oled_data = 16'b1110010011010110;
				18'b000101110000001110: oled_data = 16'b1101110011010110;
				18'b000101110010001110: oled_data = 16'b1101010010010100;
				18'b000101110100001110: oled_data = 16'b1011001101110000;
				18'b000101110110001110: oled_data = 16'b1100110000010011;
				18'b000101111000001110: oled_data = 16'b1110010011010110;
				18'b000101111010001110: oled_data = 16'b1101110011010101;
				18'b000101111100001110: oled_data = 16'b1101110011010101;
				18'b000101111110001110: oled_data = 16'b1101110011010110;
				18'b000110000000001110: oled_data = 16'b1101110011010101;
				18'b000110000010001110: oled_data = 16'b1101010001110100;
				18'b000110000100001110: oled_data = 16'b1101110011010110;
				18'b000110000110001110: oled_data = 16'b1101110011010101;
				18'b000110001000001110: oled_data = 16'b1101010010010100;
				18'b000110001010001110: oled_data = 16'b1101110011010101;
				18'b000110001100001110: oled_data = 16'b1011110100010101;
				18'b000110001110001110: oled_data = 16'b0011000110000111;
				18'b000110010000001110: oled_data = 16'b0010000101000101;
				18'b000110010010001110: oled_data = 16'b0010000100100101;
				18'b000110010100001110: oled_data = 16'b0110001010001010;
				18'b000110010110001110: oled_data = 16'b1101010010110010;
				18'b000110011000001110: oled_data = 16'b1110110100010100;
				18'b000110011010001110: oled_data = 16'b1101001111001111;
				18'b000110011100001110: oled_data = 16'b1011001010001010;
				18'b000110011110001110: oled_data = 16'b1011001000101000;
				18'b000110100000001110: oled_data = 16'b1011001000101001;
				18'b000110100010001110: oled_data = 16'b1011001000101001;
				18'b000110100100001110: oled_data = 16'b1011001000101000;
				18'b000110100110001110: oled_data = 16'b1010101000101000;
				18'b000100011000001111: oled_data = 16'b1010110000101011;
				18'b000100011010001111: oled_data = 16'b1010110000101011;
				18'b000100011100001111: oled_data = 16'b1010010000001011;
				18'b000100011110001111: oled_data = 16'b1001101110101010;
				18'b000100100000001111: oled_data = 16'b1000001101001001;
				18'b000100100010001111: oled_data = 16'b0111101011101001;
				18'b000100100100001111: oled_data = 16'b1100010100110100;
				18'b000100100110001111: oled_data = 16'b1110010100110110;
				18'b000100101000001111: oled_data = 16'b1101110011010101;
				18'b000100101010001111: oled_data = 16'b1101010010010100;
				18'b000100101100001111: oled_data = 16'b1101110011010101;
				18'b000100101110001111: oled_data = 16'b1101110011010101;
				18'b000100110000001111: oled_data = 16'b1101110011010101;
				18'b000100110010001111: oled_data = 16'b1101110011010101;
				18'b000100110100001111: oled_data = 16'b1101110010110101;
				18'b000100110110001111: oled_data = 16'b1101010001110100;
				18'b000100111000001111: oled_data = 16'b1110010011110110;
				18'b000100111010001111: oled_data = 16'b1101110011010110;
				18'b000100111100001111: oled_data = 16'b1101110011010101;
				18'b000100111110001111: oled_data = 16'b1101110011010101;
				18'b000101000000001111: oled_data = 16'b1101110011010101;
				18'b000101000010001111: oled_data = 16'b1101110010110101;
				18'b000101000100001111: oled_data = 16'b1101010001110100;
				18'b000101000110001111: oled_data = 16'b1101110011010110;
				18'b000101001000001111: oled_data = 16'b1101110011010101;
				18'b000101001010001111: oled_data = 16'b1101110010110101;
				18'b000101001100001111: oled_data = 16'b1101010001110100;
				18'b000101001110001111: oled_data = 16'b1101110011010110;
				18'b000101010000001111: oled_data = 16'b1101110011010101;
				18'b000101010010001111: oled_data = 16'b1101110011010101;
				18'b000101010100001111: oled_data = 16'b1101110011010101;
				18'b000101010110001111: oled_data = 16'b1101110011010101;
				18'b000101011000001111: oled_data = 16'b1101110011010101;
				18'b000101011010001111: oled_data = 16'b1110010011010110;
				18'b000101011100001111: oled_data = 16'b1101110011010101;
				18'b000101011110001111: oled_data = 16'b1101110011010101;
				18'b000101100000001111: oled_data = 16'b1101110011010101;
				18'b000101100010001111: oled_data = 16'b1101110011010101;
				18'b000101100100001111: oled_data = 16'b1101110011010101;
				18'b000101100110001111: oled_data = 16'b1101110011010101;
				18'b000101101000001111: oled_data = 16'b1101010011110100;
				18'b000101101010001111: oled_data = 16'b1100110011010100;
				18'b000101101100001111: oled_data = 16'b1101110010110101;
				18'b000101101110001111: oled_data = 16'b1110010011010110;
				18'b000101110000001111: oled_data = 16'b1101110011010101;
				18'b000101110010001111: oled_data = 16'b1110010011010110;
				18'b000101110100001111: oled_data = 16'b1100001111110010;
				18'b000101110110001111: oled_data = 16'b1010101101001111;
				18'b000101111000001111: oled_data = 16'b1100110000110011;
				18'b000101111010001111: oled_data = 16'b1110010011010110;
				18'b000101111100001111: oled_data = 16'b1101110011010101;
				18'b000101111110001111: oled_data = 16'b1101110011010110;
				18'b000110000000001111: oled_data = 16'b1101110011010110;
				18'b000110000010001111: oled_data = 16'b1101010010010100;
				18'b000110000100001111: oled_data = 16'b1101110010110101;
				18'b000110000110001111: oled_data = 16'b1110010011110110;
				18'b000110001000001111: oled_data = 16'b1101010010010100;
				18'b000110001010001111: oled_data = 16'b1101110010110101;
				18'b000110001100001111: oled_data = 16'b1100010011110101;
				18'b000110001110001111: oled_data = 16'b0011100111001000;
				18'b000110010000001111: oled_data = 16'b0010000100100101;
				18'b000110010010001111: oled_data = 16'b0111101100001100;
				18'b000110010100001111: oled_data = 16'b1110010100010100;
				18'b000110010110001111: oled_data = 16'b1110010010110010;
				18'b000110011000001111: oled_data = 16'b1100001100101100;
				18'b000110011010001111: oled_data = 16'b1011001001001001;
				18'b000110011100001111: oled_data = 16'b1011001000101001;
				18'b000110011110001111: oled_data = 16'b1011001000101001;
				18'b000110100000001111: oled_data = 16'b1011001000101001;
				18'b000110100010001111: oled_data = 16'b1011001000101001;
				18'b000110100100001111: oled_data = 16'b1010101000101000;
				18'b000110100110001111: oled_data = 16'b1010101000001000;
				18'b000100011000010000: oled_data = 16'b0110001011001010;
				18'b000100011010010000: oled_data = 16'b0101101010101001;
				18'b000100011100010000: oled_data = 16'b0100101001101001;
				18'b000100011110010000: oled_data = 16'b0100001000101000;
				18'b000100100000010000: oled_data = 16'b0011101000001000;
				18'b000100100010010000: oled_data = 16'b0011101000101001;
				18'b000100100100010000: oled_data = 16'b1100110100110110;
				18'b000100100110010000: oled_data = 16'b1110010011110110;
				18'b000100101000010000: oled_data = 16'b1101110011010101;
				18'b000100101010010000: oled_data = 16'b1101010010010100;
				18'b000100101100010000: oled_data = 16'b1101110011010110;
				18'b000100101110010000: oled_data = 16'b1101110011010101;
				18'b000100110000010000: oled_data = 16'b1101110011010110;
				18'b000100110010010000: oled_data = 16'b1101110011010110;
				18'b000100110100010000: oled_data = 16'b1101110010110101;
				18'b000100110110010000: oled_data = 16'b1101110010010101;
				18'b000100111000010000: oled_data = 16'b1110010011110110;
				18'b000100111010010000: oled_data = 16'b1101010010010101;
				18'b000100111100010000: oled_data = 16'b1101110010110101;
				18'b000100111110010000: oled_data = 16'b1101110011010101;
				18'b000101000000010000: oled_data = 16'b1101110011010101;
				18'b000101000010010000: oled_data = 16'b1101110010110101;
				18'b000101000100010000: oled_data = 16'b1101010001110100;
				18'b000101000110010000: oled_data = 16'b1101110011010110;
				18'b000101001000010000: oled_data = 16'b1101110011010101;
				18'b000101001010010000: oled_data = 16'b1101110011010110;
				18'b000101001100010000: oled_data = 16'b1101010001110100;
				18'b000101001110010000: oled_data = 16'b1101110011010101;
				18'b000101010000010000: oled_data = 16'b1101110011010101;
				18'b000101010010010000: oled_data = 16'b1101110011010101;
				18'b000101010100010000: oled_data = 16'b1101110011010101;
				18'b000101010110010000: oled_data = 16'b1101110011010101;
				18'b000101011000010000: oled_data = 16'b1101110011010101;
				18'b000101011010010000: oled_data = 16'b1110110101111000;
				18'b000101011100010000: oled_data = 16'b1101110011110110;
				18'b000101011110010000: oled_data = 16'b1101110011010101;
				18'b000101100000010000: oled_data = 16'b1101110011010101;
				18'b000101100010010000: oled_data = 16'b1101110011010101;
				18'b000101100100010000: oled_data = 16'b1101110010110101;
				18'b000101100110010000: oled_data = 16'b1101110011010101;
				18'b000101101000010000: oled_data = 16'b1101110011010101;
				18'b000101101010010000: oled_data = 16'b1101110111111000;
				18'b000101101100010000: oled_data = 16'b1101010100010101;
				18'b000101101110010000: oled_data = 16'b1101110011010101;
				18'b000101110000010000: oled_data = 16'b1101110011010101;
				18'b000101110010010000: oled_data = 16'b1101110011010110;
				18'b000101110100010000: oled_data = 16'b1101110010110101;
				18'b000101110110010000: oled_data = 16'b1011001101110000;
				18'b000101111000010000: oled_data = 16'b1011001101010000;
				18'b000101111010010000: oled_data = 16'b1100110001010011;
				18'b000101111100010000: oled_data = 16'b1110010011010110;
				18'b000101111110010000: oled_data = 16'b1101110011010110;
				18'b000110000000010000: oled_data = 16'b1101110011010110;
				18'b000110000010010000: oled_data = 16'b1101110010110101;
				18'b000110000100010000: oled_data = 16'b1101010010010101;
				18'b000110000110010000: oled_data = 16'b1110010011110110;
				18'b000110001000010000: oled_data = 16'b1101010010010100;
				18'b000110001010010000: oled_data = 16'b1101110010010101;
				18'b000110001100010000: oled_data = 16'b1101010011010110;
				18'b000110001110010000: oled_data = 16'b0101101001001010;
				18'b000110010000010000: oled_data = 16'b1000101100001101;
				18'b000110010010010000: oled_data = 16'b1110110100110101;
				18'b000110010100010000: oled_data = 16'b1110010001010001;
				18'b000110010110010000: oled_data = 16'b1011101010101010;
				18'b000110011000010000: oled_data = 16'b1011001000101001;
				18'b000110011010010000: oled_data = 16'b1011001001001001;
				18'b000110011100010000: oled_data = 16'b1011001000101001;
				18'b000110011110010000: oled_data = 16'b1011001000101001;
				18'b000110100000010000: oled_data = 16'b1011001000101001;
				18'b000110100010010000: oled_data = 16'b1011001000101001;
				18'b000110100100010000: oled_data = 16'b1010101000101000;
				18'b000110100110010000: oled_data = 16'b1010101000001000;
				18'b000100011000010001: oled_data = 16'b0011001001001011;
				18'b000100011010010001: oled_data = 16'b0101110001110011;
				18'b000100011100010001: oled_data = 16'b0110010100110101;
				18'b000100011110010001: oled_data = 16'b0101010001110011;
				18'b000100100000010001: oled_data = 16'b0100001101101111;
				18'b000100100010010001: oled_data = 16'b0100101011101101;
				18'b000100100100010001: oled_data = 16'b1101110100110111;
				18'b000100100110010001: oled_data = 16'b1110010011010110;
				18'b000100101000010001: oled_data = 16'b1101110010110101;
				18'b000100101010010001: oled_data = 16'b1101010010010100;
				18'b000100101100010001: oled_data = 16'b1101110011010110;
				18'b000100101110010001: oled_data = 16'b1101110011010101;
				18'b000100110000010001: oled_data = 16'b1110010011110110;
				18'b000100110010010001: oled_data = 16'b1101110011110110;
				18'b000100110100010001: oled_data = 16'b1101010010010101;
				18'b000100110110010001: oled_data = 16'b1101110010110101;
				18'b000100111000010001: oled_data = 16'b1110010011110110;
				18'b000100111010010001: oled_data = 16'b1101010001110100;
				18'b000100111100010001: oled_data = 16'b1101110010110101;
				18'b000100111110010001: oled_data = 16'b1101110011010101;
				18'b000101000000010001: oled_data = 16'b1101110011010101;
				18'b000101000010010001: oled_data = 16'b1101110010110101;
				18'b000101000100010001: oled_data = 16'b1101010001110100;
				18'b000101000110010001: oled_data = 16'b1101110011010101;
				18'b000101001000010001: oled_data = 16'b1101110011010101;
				18'b000101001010010001: oled_data = 16'b1110010011010110;
				18'b000101001100010001: oled_data = 16'b1101010010010100;
				18'b000101001110010001: oled_data = 16'b1101110010110101;
				18'b000101010000010001: oled_data = 16'b1101110011010110;
				18'b000101010010010001: oled_data = 16'b1101110011010101;
				18'b000101010100010001: oled_data = 16'b1101110011010101;
				18'b000101010110010001: oled_data = 16'b1101110011010101;
				18'b000101011000010001: oled_data = 16'b1101110010110101;
				18'b000101011010010001: oled_data = 16'b1110010101110111;
				18'b000101011100010001: oled_data = 16'b1110010101110111;
				18'b000101011110010001: oled_data = 16'b1101110011010101;
				18'b000101100000010001: oled_data = 16'b1101110011010101;
				18'b000101100010010001: oled_data = 16'b1101110011010101;
				18'b000101100100010001: oled_data = 16'b1101110010110101;
				18'b000101100110010001: oled_data = 16'b1101010001110100;
				18'b000101101000010001: oled_data = 16'b1101110011010101;
				18'b000101101010010001: oled_data = 16'b1101110101010110;
				18'b000101101100010001: oled_data = 16'b1101111010011001;
				18'b000101101110010001: oled_data = 16'b1100110100010101;
				18'b000101110000010001: oled_data = 16'b1101110011010101;
				18'b000101110010010001: oled_data = 16'b1101110011010101;
				18'b000101110100010001: oled_data = 16'b1110010011110110;
				18'b000101110110010001: oled_data = 16'b1100001111110010;
				18'b000101111000010001: oled_data = 16'b1011001101001111;
				18'b000101111010010001: oled_data = 16'b1011001101110000;
				18'b000101111100010001: oled_data = 16'b1101010010010100;
				18'b000101111110010001: oled_data = 16'b1110010011010110;
				18'b000110000000010001: oled_data = 16'b1101110011010110;
				18'b000110000010010001: oled_data = 16'b1101110011010101;
				18'b000110000100010001: oled_data = 16'b1101010001110100;
				18'b000110000110010001: oled_data = 16'b1110010011110110;
				18'b000110001000010001: oled_data = 16'b1101110010010101;
				18'b000110001010010001: oled_data = 16'b1101110010110101;
				18'b000110001100010001: oled_data = 16'b1101110010010101;
				18'b000110001110010001: oled_data = 16'b1100010000110010;
				18'b000110010000010001: oled_data = 16'b1110010100010100;
				18'b000110010010010001: oled_data = 16'b1101110000110000;
				18'b000110010100010001: oled_data = 16'b1011001010001010;
				18'b000110010110010001: oled_data = 16'b1011001000101000;
				18'b000110011000010001: oled_data = 16'b1011001001001001;
				18'b000110011010010001: oled_data = 16'b1011001000101001;
				18'b000110011100010001: oled_data = 16'b1011001000101001;
				18'b000110011110010001: oled_data = 16'b1011001000101001;
				18'b000110100000010001: oled_data = 16'b1011001000101001;
				18'b000110100010010001: oled_data = 16'b1011001000101001;
				18'b000110100100010001: oled_data = 16'b1011001000101000;
				18'b000110100110010001: oled_data = 16'b1011001000001000;
				18'b000100011000010010: oled_data = 16'b0100101101101111;
				18'b000100011010010010: oled_data = 16'b0111111000111010;
				18'b000100011100010010: oled_data = 16'b0111011001011011;
				18'b000100011110010010: oled_data = 16'b0111011000111010;
				18'b000100100000010010: oled_data = 16'b0111011000011001;
				18'b000100100010010010: oled_data = 16'b0111010111111001;
				18'b000100100100010010: oled_data = 16'b1001010110111001;
				18'b000100100110010010: oled_data = 16'b1011010100110111;
				18'b000100101000010010: oled_data = 16'b1101010010110101;
				18'b000100101010010010: oled_data = 16'b1101110010110101;
				18'b000100101100010010: oled_data = 16'b1101110011010110;
				18'b000100101110010010: oled_data = 16'b1101110011010101;
				18'b000100110000010010: oled_data = 16'b1101110011010110;
				18'b000100110010010010: oled_data = 16'b1101110011010110;
				18'b000100110100010010: oled_data = 16'b1101010010010100;
				18'b000100110110010010: oled_data = 16'b1101110010110101;
				18'b000100111000010010: oled_data = 16'b1110010011010110;
				18'b000100111010010010: oled_data = 16'b1101010001110100;
				18'b000100111100010010: oled_data = 16'b1101110011010101;
				18'b000100111110010010: oled_data = 16'b1101110011010101;
				18'b000101000000010010: oled_data = 16'b1101110011010101;
				18'b000101000010010010: oled_data = 16'b1101110011010101;
				18'b000101000100010010: oled_data = 16'b1101010001110100;
				18'b000101000110010010: oled_data = 16'b1101110011010101;
				18'b000101001000010010: oled_data = 16'b1101110011010110;
				18'b000101001010010010: oled_data = 16'b1110010011010110;
				18'b000101001100010010: oled_data = 16'b1101110010110101;
				18'b000101001110010010: oled_data = 16'b1100110001010011;
				18'b000101010000010010: oled_data = 16'b1101110011010110;
				18'b000101010010010010: oled_data = 16'b1101110011010110;
				18'b000101010100010010: oled_data = 16'b1101110011010101;
				18'b000101010110010010: oled_data = 16'b1101110011010101;
				18'b000101011000010010: oled_data = 16'b1101110011010101;
				18'b000101011010010010: oled_data = 16'b1101110011110110;
				18'b000101011100010010: oled_data = 16'b1110110110011000;
				18'b000101011110010010: oled_data = 16'b1101110011010101;
				18'b000101100000010010: oled_data = 16'b1101110011010101;
				18'b000101100010010010: oled_data = 16'b1101110011010101;
				18'b000101100100010010: oled_data = 16'b1101110011010110;
				18'b000101100110010010: oled_data = 16'b1101010010010101;
				18'b000101101000010010: oled_data = 16'b1101110010110101;
				18'b000101101010010010: oled_data = 16'b1101010011110101;
				18'b000101101100010010: oled_data = 16'b1101111010011001;
				18'b000101101110010010: oled_data = 16'b1101111010011001;
				18'b000101110000010010: oled_data = 16'b1101010011110100;
				18'b000101110010010010: oled_data = 16'b1101110011010101;
				18'b000101110100010010: oled_data = 16'b1101110011010110;
				18'b000101110110010010: oled_data = 16'b1101010010010101;
				18'b000101111000010010: oled_data = 16'b1010101101010000;
				18'b000101111010010010: oled_data = 16'b1011001101110000;
				18'b000101111100010010: oled_data = 16'b1011101110010001;
				18'b000101111110010010: oled_data = 16'b1101110010110101;
				18'b000110000000010010: oled_data = 16'b1110010011010110;
				18'b000110000010010010: oled_data = 16'b1101110011010110;
				18'b000110000100010010: oled_data = 16'b1101010001110100;
				18'b000110000110010010: oled_data = 16'b1101110011010101;
				18'b000110001000010010: oled_data = 16'b1101110010110101;
				18'b000110001010010010: oled_data = 16'b1101010010010100;
				18'b000110001100010010: oled_data = 16'b1101010001110011;
				18'b000110001110010010: oled_data = 16'b1110010011110101;
				18'b000110010000010010: oled_data = 16'b1101010000110000;
				18'b000110010010010010: oled_data = 16'b1011001001101010;
				18'b000110010100010010: oled_data = 16'b1011101001001001;
				18'b000110010110010010: oled_data = 16'b1011001001001001;
				18'b000110011000010010: oled_data = 16'b1011001001001001;
				18'b000110011010010010: oled_data = 16'b1011001001001001;
				18'b000110011100010010: oled_data = 16'b1011001000101001;
				18'b000110011110010010: oled_data = 16'b1011001000101001;
				18'b000110100000010010: oled_data = 16'b1011001000101001;
				18'b000110100010010010: oled_data = 16'b1011001000101001;
				18'b000110100100010010: oled_data = 16'b1011001000101000;
				18'b000110100110010010: oled_data = 16'b1011001000101000;
				18'b000100011000010011: oled_data = 16'b0101110001110010;
				18'b000100011010010011: oled_data = 16'b0111011000111010;
				18'b000100011100010011: oled_data = 16'b0110110111011010;
				18'b000100011110010011: oled_data = 16'b0111010111011001;
				18'b000100100000010011: oled_data = 16'b1001111010111100;
				18'b000100100010010011: oled_data = 16'b1010011011111100;
				18'b000100100100010011: oled_data = 16'b1000011001111011;
				18'b000100100110010011: oled_data = 16'b0111011000011001;
				18'b000100101000010011: oled_data = 16'b1001110101111000;
				18'b000100101010010011: oled_data = 16'b1101110011010110;
				18'b000100101100010011: oled_data = 16'b1101110011010101;
				18'b000100101110010011: oled_data = 16'b1101110011010101;
				18'b000100110000010011: oled_data = 16'b1101110011010101;
				18'b000100110010010011: oled_data = 16'b1110010011010110;
				18'b000100110100010011: oled_data = 16'b1101010001110100;
				18'b000100110110010011: oled_data = 16'b1101110010110101;
				18'b000100111000010011: oled_data = 16'b1101110011010110;
				18'b000100111010010011: oled_data = 16'b1101010001110100;
				18'b000100111100010011: oled_data = 16'b1101110011010101;
				18'b000100111110010011: oled_data = 16'b1101110011010101;
				18'b000101000000010011: oled_data = 16'b1101110011010101;
				18'b000101000010010011: oled_data = 16'b1101110011010110;
				18'b000101000100010011: oled_data = 16'b1101010001110100;
				18'b000101000110010011: oled_data = 16'b1101110010110101;
				18'b000101001000010011: oled_data = 16'b1110010011110110;
				18'b000101001010010011: oled_data = 16'b1110010011010110;
				18'b000101001100010011: oled_data = 16'b1101110011010101;
				18'b000101001110010011: oled_data = 16'b1100010000010010;
				18'b000101010000010011: oled_data = 16'b1101110011010101;
				18'b000101010010010011: oled_data = 16'b1101110011010110;
				18'b000101010100010011: oled_data = 16'b1101110011010110;
				18'b000101010110010011: oled_data = 16'b1101110011010101;
				18'b000101011000010011: oled_data = 16'b1101110011010101;
				18'b000101011010010011: oled_data = 16'b1101110011010101;
				18'b000101011100010011: oled_data = 16'b1110010100010110;
				18'b000101011110010011: oled_data = 16'b1101110011010110;
				18'b000101100000010011: oled_data = 16'b1101110011010101;
				18'b000101100010010011: oled_data = 16'b1101110011010101;
				18'b000101100100010011: oled_data = 16'b1101110011010101;
				18'b000101100110010011: oled_data = 16'b1101110011010101;
				18'b000101101000010011: oled_data = 16'b1101010001110100;
				18'b000101101010010011: oled_data = 16'b1101110010110101;
				18'b000101101100010011: oled_data = 16'b1101110110110111;
				18'b000101101110010011: oled_data = 16'b1110111100111011;
				18'b000101110000010011: oled_data = 16'b1101111000010111;
				18'b000101110010010011: oled_data = 16'b1101010011010101;
				18'b000101110100010011: oled_data = 16'b1101110011010101;
				18'b000101110110010011: oled_data = 16'b1101110011110110;
				18'b000101111000010011: oled_data = 16'b1100110011010101;
				18'b000101111010010011: oled_data = 16'b1011001111010001;
				18'b000101111100010011: oled_data = 16'b1011101110010001;
				18'b000101111110010011: oled_data = 16'b1100001111110010;
				18'b000110000000010011: oled_data = 16'b1101110011010101;
				18'b000110000010010011: oled_data = 16'b1101110011010110;
				18'b000110000100010011: oled_data = 16'b1101010010010100;
				18'b000110000110010011: oled_data = 16'b1101110010110101;
				18'b000110001000010011: oled_data = 16'b1101010010010100;
				18'b000110001010010011: oled_data = 16'b1100110000110010;
				18'b000110001100010011: oled_data = 16'b1110010011110100;
				18'b000110001110010011: oled_data = 16'b1101110001010001;
				18'b000110010000010011: oled_data = 16'b1011101010001010;
				18'b000110010010010011: oled_data = 16'b1011001001001001;
				18'b000110010100010011: oled_data = 16'b1011101001001001;
				18'b000110010110010011: oled_data = 16'b1011001001001001;
				18'b000110011000010011: oled_data = 16'b1011001001001001;
				18'b000110011010010011: oled_data = 16'b1011001001001001;
				18'b000110011100010011: oled_data = 16'b1011001001001001;
				18'b000110011110010011: oled_data = 16'b1011001000101001;
				18'b000110100000010011: oled_data = 16'b1011001000101001;
				18'b000110100010010011: oled_data = 16'b1011001000101001;
				18'b000110100100010011: oled_data = 16'b1011001000101000;
				18'b000110100110010011: oled_data = 16'b1011001000101000;
				18'b000100011000010100: oled_data = 16'b0110010100010101;
				18'b000100011010010100: oled_data = 16'b0111011000011010;
				18'b000100011100010100: oled_data = 16'b0101010011110111;
				18'b000100011110010100: oled_data = 16'b1000111001011010;
				18'b000100100000010100: oled_data = 16'b1011111100111101;
				18'b000100100010010100: oled_data = 16'b1001011000011010;
				18'b000100100100010100: oled_data = 16'b0101110010110110;
				18'b000100100110010100: oled_data = 16'b0111010111111010;
				18'b000100101000010100: oled_data = 16'b0111111000011001;
				18'b000100101010010100: oled_data = 16'b1101010011110110;
				18'b000100101100010100: oled_data = 16'b1101110011010101;
				18'b000100101110010100: oled_data = 16'b1101110011010101;
				18'b000100110000010100: oled_data = 16'b1101110011010101;
				18'b000100110010010100: oled_data = 16'b1110010011010110;
				18'b000100110100010100: oled_data = 16'b1101010010010100;
				18'b000100110110010100: oled_data = 16'b1101110010110101;
				18'b000100111000010100: oled_data = 16'b1101110011010101;
				18'b000100111010010100: oled_data = 16'b1101010001010100;
				18'b000100111100010100: oled_data = 16'b1101110011010101;
				18'b000100111110010100: oled_data = 16'b1101110011010101;
				18'b000101000000010100: oled_data = 16'b1101110011010101;
				18'b000101000010010100: oled_data = 16'b1101110011010110;
				18'b000101000100010100: oled_data = 16'b1101110010010101;
				18'b000101000110010100: oled_data = 16'b1101110010010101;
				18'b000101001000010100: oled_data = 16'b1110010011010110;
				18'b000101001010010100: oled_data = 16'b1110010011010110;
				18'b000101001100010100: oled_data = 16'b1101110011010110;
				18'b000101001110010100: oled_data = 16'b1100110001110100;
				18'b000101010000010100: oled_data = 16'b1101010010010100;
				18'b000101010010010100: oled_data = 16'b1101110011010110;
				18'b000101010100010100: oled_data = 16'b1101110011010101;
				18'b000101010110010100: oled_data = 16'b1101110011010101;
				18'b000101011000010100: oled_data = 16'b1101110011010101;
				18'b000101011010010100: oled_data = 16'b1101110011010101;
				18'b000101011100010100: oled_data = 16'b1101110011010101;
				18'b000101011110010100: oled_data = 16'b1101110011010101;
				18'b000101100000010100: oled_data = 16'b1101110011010101;
				18'b000101100010010100: oled_data = 16'b1101110011010101;
				18'b000101100100010100: oled_data = 16'b1101110011010101;
				18'b000101100110010100: oled_data = 16'b1101110011010110;
				18'b000101101000010100: oled_data = 16'b1101010010010101;
				18'b000101101010010100: oled_data = 16'b1101010001110100;
				18'b000101101100010100: oled_data = 16'b1101010100110101;
				18'b000101101110010100: oled_data = 16'b1110111011111010;
				18'b000101110000010100: oled_data = 16'b1110111100011011;
				18'b000101110010010100: oled_data = 16'b1101010101110110;
				18'b000101110100010100: oled_data = 16'b1101110011010101;
				18'b000101110110010100: oled_data = 16'b1101110011010110;
				18'b000101111000010100: oled_data = 16'b1101010100110110;
				18'b000101111010010100: oled_data = 16'b1100110101110110;
				18'b000101111100010100: oled_data = 16'b1011001110010000;
				18'b000101111110010100: oled_data = 16'b1011001110010001;
				18'b000110000000010100: oled_data = 16'b1100110000010011;
				18'b000110000010010100: oled_data = 16'b1110010011010110;
				18'b000110000100010100: oled_data = 16'b1101110010010101;
				18'b000110000110010100: oled_data = 16'b1101010010010100;
				18'b000110001000010100: oled_data = 16'b1101010001110011;
				18'b000110001010010100: oled_data = 16'b1110010011010100;
				18'b000110001100010100: oled_data = 16'b1110110010110011;
				18'b000110001110010100: oled_data = 16'b1011101010101011;
				18'b000110010000010100: oled_data = 16'b1011001001001001;
				18'b000110010010010100: oled_data = 16'b1011101001001001;
				18'b000110010100010100: oled_data = 16'b1011001001001001;
				18'b000110010110010100: oled_data = 16'b1011001001001001;
				18'b000110011000010100: oled_data = 16'b1011001001001001;
				18'b000110011010010100: oled_data = 16'b1011001001001001;
				18'b000110011100010100: oled_data = 16'b1011001001001001;
				18'b000110011110010100: oled_data = 16'b1011001000101001;
				18'b000110100000010100: oled_data = 16'b1011001000101000;
				18'b000110100010010100: oled_data = 16'b1011001000101001;
				18'b000110100100010100: oled_data = 16'b1011001000101000;
				18'b000110100110010100: oled_data = 16'b1011001000101000;
				18'b000100011000010101: oled_data = 16'b0110110110110111;
				18'b000100011010010101: oled_data = 16'b0110010101111000;
				18'b000100011100010101: oled_data = 16'b0100110010010110;
				18'b000100011110010101: oled_data = 16'b1010011010111011;
				18'b000100100000010101: oled_data = 16'b1010111010111011;
				18'b000100100010010101: oled_data = 16'b0101010010010110;
				18'b000100100100010101: oled_data = 16'b0100010001010101;
				18'b000100100110010101: oled_data = 16'b0101110100110111;
				18'b000100101000010101: oled_data = 16'b1000010111111001;
				18'b000100101010010101: oled_data = 16'b1101010011010110;
				18'b000100101100010101: oled_data = 16'b1101110011010101;
				18'b000100101110010101: oled_data = 16'b1101110011010101;
				18'b000100110000010101: oled_data = 16'b1101110011010101;
				18'b000100110010010101: oled_data = 16'b1101110011010110;
				18'b000100110100010101: oled_data = 16'b1101010001110100;
				18'b000100110110010101: oled_data = 16'b1101110010110101;
				18'b000100111000010101: oled_data = 16'b1101110011010101;
				18'b000100111010010101: oled_data = 16'b1100110000110011;
				18'b000100111100010101: oled_data = 16'b1101110011010101;
				18'b000100111110010101: oled_data = 16'b1101110011010101;
				18'b000101000000010101: oled_data = 16'b1101110011010101;
				18'b000101000010010101: oled_data = 16'b1101110011010101;
				18'b000101000100010101: oled_data = 16'b1101110010110101;
				18'b000101000110010101: oled_data = 16'b1101010010010100;
				18'b000101001000010101: oled_data = 16'b1101110011010110;
				18'b000101001010010101: oled_data = 16'b1101110011010110;
				18'b000101001100010101: oled_data = 16'b1101110011010110;
				18'b000101001110010101: oled_data = 16'b1101010010110101;
				18'b000101010000010101: oled_data = 16'b1100010001010011;
				18'b000101010010010101: oled_data = 16'b1101110011010101;
				18'b000101010100010101: oled_data = 16'b1101110011010101;
				18'b000101010110010101: oled_data = 16'b1101110011010101;
				18'b000101011000010101: oled_data = 16'b1101110011010101;
				18'b000101011010010101: oled_data = 16'b1101110011010101;
				18'b000101011100010101: oled_data = 16'b1101110011010101;
				18'b000101011110010101: oled_data = 16'b1101110011010101;
				18'b000101100000010101: oled_data = 16'b1101110011010101;
				18'b000101100010010101: oled_data = 16'b1101110011010101;
				18'b000101100100010101: oled_data = 16'b1101110011010101;
				18'b000101100110010101: oled_data = 16'b1101110011010101;
				18'b000101101000010101: oled_data = 16'b1101110011010101;
				18'b000101101010010101: oled_data = 16'b1101010001110100;
				18'b000101101100010101: oled_data = 16'b1101010010110100;
				18'b000101101110010101: oled_data = 16'b1110011010011010;
				18'b000101110000010101: oled_data = 16'b1110011011011010;
				18'b000101110010010101: oled_data = 16'b1101011001011000;
				18'b000101110100010101: oled_data = 16'b1100110011110100;
				18'b000101110110010101: oled_data = 16'b1101110011010110;
				18'b000101111000010101: oled_data = 16'b1101010011110101;
				18'b000101111010010101: oled_data = 16'b1101111000011000;
				18'b000101111100010101: oled_data = 16'b1010101110010000;
				18'b000101111110010101: oled_data = 16'b1011001110010001;
				18'b000110000000010101: oled_data = 16'b1011001110010001;
				18'b000110000010010101: oled_data = 16'b1101010001110101;
				18'b000110000100010101: oled_data = 16'b1101110010110101;
				18'b000110000110010101: oled_data = 16'b1011001110110000;
				18'b000110001000010101: oled_data = 16'b1101110010110011;
				18'b000110001010010101: oled_data = 16'b1110110100010100;
				18'b000110001100010101: oled_data = 16'b1100001100101101;
				18'b000110001110010101: oled_data = 16'b1011001000101001;
				18'b000110010000010101: oled_data = 16'b1011001001001001;
				18'b000110010010010101: oled_data = 16'b1011001001001001;
				18'b000110010100010101: oled_data = 16'b1011001001001001;
				18'b000110010110010101: oled_data = 16'b1011001001001001;
				18'b000110011000010101: oled_data = 16'b1011001001001001;
				18'b000110011010010101: oled_data = 16'b1011001001001001;
				18'b000110011100010101: oled_data = 16'b1011001000101001;
				18'b000110011110010101: oled_data = 16'b1010001000001000;
				18'b000110100000010101: oled_data = 16'b1010101000101000;
				18'b000110100010010101: oled_data = 16'b1011001000101001;
				18'b000110100100010101: oled_data = 16'b1011001000101000;
				18'b000110100110010101: oled_data = 16'b1011001000101000;
				18'b000100011000010110: oled_data = 16'b0111010111111001;
				18'b000100011010010110: oled_data = 16'b0101010011110111;
				18'b000100011100010110: oled_data = 16'b0100110010010110;
				18'b000100011110010110: oled_data = 16'b1001111010011100;
				18'b000100100000010110: oled_data = 16'b0111110101010111;
				18'b000100100010010110: oled_data = 16'b0100110001010101;
				18'b000100100100010110: oled_data = 16'b0100110001010110;
				18'b000100100110010110: oled_data = 16'b0101010011010110;
				18'b000100101000010110: oled_data = 16'b1000010111011001;
				18'b000100101010010110: oled_data = 16'b1101010011010101;
				18'b000100101100010110: oled_data = 16'b1101110011010101;
				18'b000100101110010110: oled_data = 16'b1101110011010101;
				18'b000100110000010110: oled_data = 16'b1101110011010101;
				18'b000100110010010110: oled_data = 16'b1101110011010110;
				18'b000100110100010110: oled_data = 16'b1101010001110100;
				18'b000100110110010110: oled_data = 16'b1101110010110101;
				18'b000100111000010110: oled_data = 16'b1101110011010101;
				18'b000100111010010110: oled_data = 16'b1100110000110011;
				18'b000100111100010110: oled_data = 16'b1101110011010101;
				18'b000100111110010110: oled_data = 16'b1101110011010101;
				18'b000101000000010110: oled_data = 16'b1101110011010101;
				18'b000101000010010110: oled_data = 16'b1101110011010101;
				18'b000101000100010110: oled_data = 16'b1101110011010110;
				18'b000101000110010110: oled_data = 16'b1100110000110011;
				18'b000101001000010110: oled_data = 16'b1101110010110101;
				18'b000101001010010110: oled_data = 16'b1101110011010101;
				18'b000101001100010110: oled_data = 16'b1101110011010101;
				18'b000101001110010110: oled_data = 16'b1101110011010101;
				18'b000101010000010110: oled_data = 16'b1100110001110011;
				18'b000101010010010110: oled_data = 16'b1101010010110101;
				18'b000101010100010110: oled_data = 16'b1101110011010101;
				18'b000101010110010110: oled_data = 16'b1101110011010101;
				18'b000101011000010110: oled_data = 16'b1101110011010101;
				18'b000101011010010110: oled_data = 16'b1101110011010101;
				18'b000101011100010110: oled_data = 16'b1101110011010101;
				18'b000101011110010110: oled_data = 16'b1101110011010101;
				18'b000101100000010110: oled_data = 16'b1101110011010101;
				18'b000101100010010110: oled_data = 16'b1101110011010101;
				18'b000101100100010110: oled_data = 16'b1101110011010101;
				18'b000101100110010110: oled_data = 16'b1101110011010110;
				18'b000101101000010110: oled_data = 16'b1110010011010110;
				18'b000101101010010110: oled_data = 16'b1101010010010100;
				18'b000101101100010110: oled_data = 16'b1101010001110100;
				18'b000101101110010110: oled_data = 16'b1101010110010110;
				18'b000101110000010110: oled_data = 16'b1101111010111001;
				18'b000101110010010110: oled_data = 16'b1110011011111010;
				18'b000101110100010110: oled_data = 16'b1010010001010001;
				18'b000101110110010110: oled_data = 16'b1101010010110101;
				18'b000101111000010110: oled_data = 16'b1101110011010101;
				18'b000101111010010110: oled_data = 16'b1101010111010111;
				18'b000101111100010110: oled_data = 16'b1011010000110010;
				18'b000101111110010110: oled_data = 16'b1010101100110000;
				18'b000110000000010110: oled_data = 16'b1011101110010001;
				18'b000110000010010110: oled_data = 16'b1011101111010010;
				18'b000110000100010110: oled_data = 16'b1101110010110101;
				18'b000110000110010110: oled_data = 16'b1011101111110001;
				18'b000110001000010110: oled_data = 16'b1110110100010100;
				18'b000110001010010110: oled_data = 16'b1101001111101111;
				18'b000110001100010110: oled_data = 16'b1011001001001001;
				18'b000110001110010110: oled_data = 16'b1011001001001001;
				18'b000110010000010110: oled_data = 16'b1011001001001001;
				18'b000110010010010110: oled_data = 16'b1011001001001001;
				18'b000110010100010110: oled_data = 16'b1011001001001001;
				18'b000110010110010110: oled_data = 16'b1011001001001001;
				18'b000110011000010110: oled_data = 16'b1011001001001001;
				18'b000110011010010110: oled_data = 16'b1011001000101001;
				18'b000110011100010110: oled_data = 16'b1010100111101000;
				18'b000110011110010110: oled_data = 16'b1011001000101000;
				18'b000110100000010110: oled_data = 16'b1011001000101001;
				18'b000110100010010110: oled_data = 16'b1011001000101001;
				18'b000110100100010110: oled_data = 16'b1011001000101000;
				18'b000110100110010110: oled_data = 16'b1011001000101000;
				18'b000100011000010111: oled_data = 16'b0111011000011001;
				18'b000100011010010111: oled_data = 16'b0101010010110110;
				18'b000100011100010111: oled_data = 16'b0100110001010101;
				18'b000100011110010111: oled_data = 16'b0110110100111000;
				18'b000100100000010111: oled_data = 16'b0101010001110110;
				18'b000100100010010111: oled_data = 16'b0100110001010101;
				18'b000100100100010111: oled_data = 16'b0100110001010101;
				18'b000100100110010111: oled_data = 16'b0101010010110110;
				18'b000100101000010111: oled_data = 16'b1000110110011000;
				18'b000100101010010111: oled_data = 16'b1101110011010101;
				18'b000100101100010111: oled_data = 16'b1101110011010101;
				18'b000100101110010111: oled_data = 16'b1101110011010101;
				18'b000100110000010111: oled_data = 16'b1101110011010101;
				18'b000100110010010111: oled_data = 16'b1101110011010110;
				18'b000100110100010111: oled_data = 16'b1101010001110100;
				18'b000100110110010111: oled_data = 16'b1101110010110101;
				18'b000100111000010111: oled_data = 16'b1101110011010101;
				18'b000100111010010111: oled_data = 16'b1100110000110011;
				18'b000100111100010111: oled_data = 16'b1101110010110101;
				18'b000100111110010111: oled_data = 16'b1101110011010101;
				18'b000101000000010111: oled_data = 16'b1101110011010101;
				18'b000101000010010111: oled_data = 16'b1101110011010101;
				18'b000101000100010111: oled_data = 16'b1110010011010110;
				18'b000101000110010111: oled_data = 16'b1100110001110100;
				18'b000101001000010111: oled_data = 16'b1101010010010100;
				18'b000101001010010111: oled_data = 16'b1110010011010110;
				18'b000101001100010111: oled_data = 16'b1101110011010101;
				18'b000101001110010111: oled_data = 16'b1101110011010101;
				18'b000101010000010111: oled_data = 16'b1101010011010101;
				18'b000101010010010111: oled_data = 16'b1100110011110101;
				18'b000101010100010111: oled_data = 16'b1101110010110101;
				18'b000101010110010111: oled_data = 16'b1101110011010101;
				18'b000101011000010111: oled_data = 16'b1101110011010101;
				18'b000101011010010111: oled_data = 16'b1101110011010101;
				18'b000101011100010111: oled_data = 16'b1101110011010101;
				18'b000101011110010111: oled_data = 16'b1101110011010101;
				18'b000101100000010111: oled_data = 16'b1101110011010101;
				18'b000101100010010111: oled_data = 16'b1101110011010101;
				18'b000101100100010111: oled_data = 16'b1101110011010101;
				18'b000101100110010111: oled_data = 16'b1101110010010101;
				18'b000101101000010111: oled_data = 16'b1101010001110100;
				18'b000101101010010111: oled_data = 16'b1100110001010011;
				18'b000101101100010111: oled_data = 16'b1100010000010011;
				18'b000101101110010111: oled_data = 16'b1101010110010111;
				18'b000101110000010111: oled_data = 16'b1110111101011011;
				18'b000101110010010111: oled_data = 16'b1100111000010111;
				18'b000101110100010111: oled_data = 16'b0110001011001010;
				18'b000101110110010111: oled_data = 16'b1100110011110101;
				18'b000101111000010111: oled_data = 16'b1101110011010110;
				18'b000101111010010111: oled_data = 16'b1101010101110111;
				18'b000101111100010111: oled_data = 16'b1100010011010100;
				18'b000101111110010111: oled_data = 16'b1010101100110000;
				18'b000110000000010111: oled_data = 16'b1011001101110001;
				18'b000110000010010111: oled_data = 16'b1011101110010001;
				18'b000110000100010111: oled_data = 16'b1100010000010010;
				18'b000110000110010111: oled_data = 16'b1110010011110100;
				18'b000110001000010111: oled_data = 16'b1110010010110010;
				18'b000110001010010111: oled_data = 16'b1011101010001010;
				18'b000110001100010111: oled_data = 16'b1011001001001001;
				18'b000110001110010111: oled_data = 16'b1011101001001001;
				18'b000110010000010111: oled_data = 16'b1011001001001001;
				18'b000110010010010111: oled_data = 16'b1011001001001001;
				18'b000110010100010111: oled_data = 16'b1011001001001001;
				18'b000110010110010111: oled_data = 16'b1011001001001001;
				18'b000110011000010111: oled_data = 16'b1011001000101001;
				18'b000110011010010111: oled_data = 16'b1010101000001000;
				18'b000110011100010111: oled_data = 16'b1011001000101001;
				18'b000110011110010111: oled_data = 16'b1011001000101001;
				18'b000110100000010111: oled_data = 16'b1011001000101001;
				18'b000110100010010111: oled_data = 16'b1011001000101000;
				18'b000110100100010111: oled_data = 16'b1011001000101000;
				18'b000110100110010111: oled_data = 16'b1010101000101000;
				18'b000100011000011000: oled_data = 16'b0111011000011010;
				18'b000100011010011000: oled_data = 16'b0101010010110110;
				18'b000100011100011000: oled_data = 16'b0100110001010110;
				18'b000100011110011000: oled_data = 16'b0100110001010110;
				18'b000100100000011000: oled_data = 16'b0100110001110110;
				18'b000100100010011000: oled_data = 16'b0100110001010110;
				18'b000100100100011000: oled_data = 16'b0100010001010101;
				18'b000100100110011000: oled_data = 16'b0101010011110110;
				18'b000100101000011000: oled_data = 16'b1001110101111000;
				18'b000100101010011000: oled_data = 16'b1101110011010101;
				18'b000100101100011000: oled_data = 16'b1101110011010101;
				18'b000100101110011000: oled_data = 16'b1101110011010101;
				18'b000100110000011000: oled_data = 16'b1101110011010101;
				18'b000100110010011000: oled_data = 16'b1101110011010110;
				18'b000100110100011000: oled_data = 16'b1101010010010100;
				18'b000100110110011000: oled_data = 16'b1101110010110101;
				18'b000100111000011000: oled_data = 16'b1101110011010101;
				18'b000100111010011000: oled_data = 16'b1100110000110011;
				18'b000100111100011000: oled_data = 16'b1101110010110101;
				18'b000100111110011000: oled_data = 16'b1101110011010101;
				18'b000101000000011000: oled_data = 16'b1101110011010101;
				18'b000101000010011000: oled_data = 16'b1101110011010101;
				18'b000101000100011000: oled_data = 16'b1110010011010110;
				18'b000101000110011000: oled_data = 16'b1101010010110101;
				18'b000101001000011000: oled_data = 16'b1100110001110100;
				18'b000101001010011000: oled_data = 16'b1101110011010101;
				18'b000101001100011000: oled_data = 16'b1101110011010101;
				18'b000101001110011000: oled_data = 16'b1101110011010101;
				18'b000101010000011000: oled_data = 16'b1101110011010101;
				18'b000101010010011000: oled_data = 16'b1101010110110111;
				18'b000101010100011000: oled_data = 16'b1101010011010101;
				18'b000101010110011000: oled_data = 16'b1101110011010101;
				18'b000101011000011000: oled_data = 16'b1101110011010101;
				18'b000101011010011000: oled_data = 16'b1101110011010101;
				18'b000101011100011000: oled_data = 16'b1101110011010101;
				18'b000101011110011000: oled_data = 16'b1101110011010101;
				18'b000101100000011000: oled_data = 16'b1101110011010101;
				18'b000101100010011000: oled_data = 16'b1101110011010101;
				18'b000101100100011000: oled_data = 16'b1101110011010101;
				18'b000101100110011000: oled_data = 16'b1101110010110101;
				18'b000101101000011000: oled_data = 16'b1101110010110101;
				18'b000101101010011000: oled_data = 16'b1101110011010101;
				18'b000101101100011000: oled_data = 16'b1101010010010100;
				18'b000101101110011000: oled_data = 16'b1101010101110110;
				18'b000101110000011000: oled_data = 16'b1110111101011011;
				18'b000101110010011000: oled_data = 16'b1000110000001111;
				18'b000101110100011000: oled_data = 16'b0011100110000101;
				18'b000101110110011000: oled_data = 16'b1011110101110101;
				18'b000101111000011000: oled_data = 16'b1101010100010101;
				18'b000101111010011000: oled_data = 16'b1101110101010110;
				18'b000101111100011000: oled_data = 16'b1100110101010110;
				18'b000101111110011000: oled_data = 16'b1011001101110000;
				18'b000110000000011000: oled_data = 16'b1011001101010000;
				18'b000110000010011000: oled_data = 16'b1011001101110001;
				18'b000110000100011000: oled_data = 16'b1100110001010010;
				18'b000110000110011000: oled_data = 16'b1110010100010100;
				18'b000110001000011000: oled_data = 16'b1100101101001101;
				18'b000110001010011000: oled_data = 16'b1011001000101000;
				18'b000110001100011000: oled_data = 16'b1011001001001001;
				18'b000110001110011000: oled_data = 16'b1011001001001001;
				18'b000110010000011000: oled_data = 16'b1011001001001001;
				18'b000110010010011000: oled_data = 16'b1011001001001001;
				18'b000110010100011000: oled_data = 16'b1011001001001001;
				18'b000110010110011000: oled_data = 16'b1011001000101001;
				18'b000110011000011000: oled_data = 16'b1010101000001000;
				18'b000110011010011000: oled_data = 16'b1011001000101001;
				18'b000110011100011000: oled_data = 16'b1011001000101001;
				18'b000110011110011000: oled_data = 16'b1011001000101001;
				18'b000110100000011000: oled_data = 16'b1011001000101001;
				18'b000110100010011000: oled_data = 16'b1011001000101000;
				18'b000110100100011000: oled_data = 16'b1011001000101000;
				18'b000110100110011000: oled_data = 16'b1010101000101000;
				18'b000100011000011001: oled_data = 16'b0111011000011010;
				18'b000100011010011001: oled_data = 16'b0101010011110111;
				18'b000100011100011001: oled_data = 16'b0100010001010110;
				18'b000100011110011001: oled_data = 16'b0100010001110110;
				18'b000100100000011001: oled_data = 16'b0100010001110110;
				18'b000100100010011001: oled_data = 16'b0100010001110110;
				18'b000100100100011001: oled_data = 16'b0100010001010101;
				18'b000100100110011001: oled_data = 16'b0110010101111000;
				18'b000100101000011001: oled_data = 16'b1010010101010111;
				18'b000100101010011001: oled_data = 16'b1110010011010101;
				18'b000100101100011001: oled_data = 16'b1101110011010110;
				18'b000100101110011001: oled_data = 16'b1101110011010101;
				18'b000100110000011001: oled_data = 16'b1101110011010101;
				18'b000100110010011001: oled_data = 16'b1101110011010110;
				18'b000100110100011001: oled_data = 16'b1101010010010100;
				18'b000100110110011001: oled_data = 16'b1101110010110101;
				18'b000100111000011001: oled_data = 16'b1101110011010110;
				18'b000100111010011001: oled_data = 16'b1100110000110011;
				18'b000100111100011001: oled_data = 16'b1101110010110101;
				18'b000100111110011001: oled_data = 16'b1101110011010110;
				18'b000101000000011001: oled_data = 16'b1101110011010101;
				18'b000101000010011001: oled_data = 16'b1101110011010101;
				18'b000101000100011001: oled_data = 16'b1101110011010101;
				18'b000101000110011001: oled_data = 16'b1101110010110101;
				18'b000101001000011001: oled_data = 16'b1101010100010101;
				18'b000101001010011001: oled_data = 16'b1101010010010100;
				18'b000101001100011001: oled_data = 16'b1110010011010110;
				18'b000101001110011001: oled_data = 16'b1101110011010101;
				18'b000101010000011001: oled_data = 16'b1101110010110101;
				18'b000101010010011001: oled_data = 16'b1101010101110110;
				18'b000101010100011001: oled_data = 16'b1101111000011000;
				18'b000101010110011001: oled_data = 16'b1101010010110100;
				18'b000101011000011001: oled_data = 16'b1101110011010101;
				18'b000101011010011001: oled_data = 16'b1101110011010101;
				18'b000101011100011001: oled_data = 16'b1101110011010101;
				18'b000101011110011001: oled_data = 16'b1101110011010101;
				18'b000101100000011001: oled_data = 16'b1101110011010101;
				18'b000101100010011001: oled_data = 16'b1101110011010101;
				18'b000101100100011001: oled_data = 16'b1101110011010101;
				18'b000101100110011001: oled_data = 16'b1101110011010101;
				18'b000101101000011001: oled_data = 16'b1101110011010101;
				18'b000101101010011001: oled_data = 16'b1101110011010110;
				18'b000101101100011001: oled_data = 16'b1101010010010100;
				18'b000101101110011001: oled_data = 16'b1100110100110101;
				18'b000101110000011001: oled_data = 16'b1101111010111001;
				18'b000101110010011001: oled_data = 16'b0101001000101000;
				18'b000101110100011001: oled_data = 16'b0101001001001000;
				18'b000101110110011001: oled_data = 16'b1101111011011001;
				18'b000101111000011001: oled_data = 16'b1101010111010111;
				18'b000101111010011001: oled_data = 16'b1101010100010101;
				18'b000101111100011001: oled_data = 16'b1101010111010111;
				18'b000101111110011001: oled_data = 16'b1011001110010001;
				18'b000110000000011001: oled_data = 16'b1011001101010000;
				18'b000110000010011001: oled_data = 16'b1011101110110001;
				18'b000110000100011001: oled_data = 16'b1110010100010100;
				18'b000110000110011001: oled_data = 16'b1101110001010001;
				18'b000110001000011001: oled_data = 16'b1011101001101010;
				18'b000110001010011001: oled_data = 16'b1011001001001001;
				18'b000110001100011001: oled_data = 16'b1011001001001001;
				18'b000110001110011001: oled_data = 16'b1011001001001001;
				18'b000110010000011001: oled_data = 16'b1011001001001001;
				18'b000110010010011001: oled_data = 16'b1011001001001001;
				18'b000110010100011001: oled_data = 16'b1011001001001001;
				18'b000110010110011001: oled_data = 16'b1010101000001000;
				18'b000110011000011001: oled_data = 16'b1011001000101001;
				18'b000110011010011001: oled_data = 16'b1011001000101001;
				18'b000110011100011001: oled_data = 16'b1011001000101001;
				18'b000110011110011001: oled_data = 16'b1011001000101000;
				18'b000110100000011001: oled_data = 16'b1011001000101001;
				18'b000110100010011001: oled_data = 16'b1011001000101000;
				18'b000110100100011001: oled_data = 16'b1011001000101000;
				18'b000110100110011001: oled_data = 16'b1010101000101000;
				18'b000100011000011010: oled_data = 16'b0111111000011010;
				18'b000100011010011010: oled_data = 16'b0110110110111001;
				18'b000100011100011010: oled_data = 16'b0100010001110101;
				18'b000100011110011010: oled_data = 16'b0100010001110101;
				18'b000100100000011010: oled_data = 16'b0100010001110101;
				18'b000100100010011010: oled_data = 16'b0100010001010110;
				18'b000100100100011010: oled_data = 16'b0100110010010110;
				18'b000100100110011010: oled_data = 16'b0110110111111010;
				18'b000100101000011010: oled_data = 16'b1010010100010110;
				18'b000100101010011010: oled_data = 16'b1110010011010101;
				18'b000100101100011010: oled_data = 16'b1101110011010110;
				18'b000100101110011010: oled_data = 16'b1101110011010101;
				18'b000100110000011010: oled_data = 16'b1101110011010101;
				18'b000100110010011010: oled_data = 16'b1101110011010110;
				18'b000100110100011010: oled_data = 16'b1101010010010100;
				18'b000100110110011010: oled_data = 16'b1101110010110101;
				18'b000100111000011010: oled_data = 16'b1101110011010110;
				18'b000100111010011010: oled_data = 16'b1101010001010100;
				18'b000100111100011010: oled_data = 16'b1101010010010101;
				18'b000100111110011010: oled_data = 16'b1101110011010110;
				18'b000101000000011010: oled_data = 16'b1101110011010101;
				18'b000101000010011010: oled_data = 16'b1101110011010101;
				18'b000101000100011010: oled_data = 16'b1101110011010101;
				18'b000101000110011010: oled_data = 16'b1101110010110101;
				18'b000101001000011010: oled_data = 16'b1110010111011000;
				18'b000101001010011010: oled_data = 16'b1100110100010101;
				18'b000101001100011010: oled_data = 16'b1101110010110101;
				18'b000101001110011010: oled_data = 16'b1101110011010101;
				18'b000101010000011010: oled_data = 16'b1101110011010101;
				18'b000101010010011010: oled_data = 16'b1101010010110101;
				18'b000101010100011010: oled_data = 16'b1110011001111010;
				18'b000101010110011010: oled_data = 16'b1101010111010111;
				18'b000101011000011010: oled_data = 16'b1101010010110101;
				18'b000101011010011010: oled_data = 16'b1101010010010101;
				18'b000101011100011010: oled_data = 16'b1101110011010101;
				18'b000101011110011010: oled_data = 16'b1101110011010101;
				18'b000101100000011010: oled_data = 16'b1101110011010101;
				18'b000101100010011010: oled_data = 16'b1101110011010101;
				18'b000101100100011010: oled_data = 16'b1101110011010101;
				18'b000101100110011010: oled_data = 16'b1101110011010101;
				18'b000101101000011010: oled_data = 16'b1101110011010101;
				18'b000101101010011010: oled_data = 16'b1101110011010110;
				18'b000101101100011010: oled_data = 16'b1101010010010100;
				18'b000101101110011010: oled_data = 16'b1100110100010101;
				18'b000101110000011010: oled_data = 16'b1010110100010011;
				18'b000101110010011010: oled_data = 16'b0011000101000101;
				18'b000101110100011010: oled_data = 16'b1001110010010001;
				18'b000101110110011010: oled_data = 16'b1110111100111011;
				18'b000101111000011010: oled_data = 16'b1110011010111001;
				18'b000101111010011010: oled_data = 16'b1100110100110101;
				18'b000101111100011010: oled_data = 16'b1101111001111001;
				18'b000101111110011010: oled_data = 16'b1011001111110010;
				18'b000110000000011010: oled_data = 16'b1011001101110000;
				18'b000110000010011010: oled_data = 16'b1101010010010010;
				18'b000110000100011010: oled_data = 16'b1110110011110100;
				18'b000110000110011010: oled_data = 16'b1100001100101101;
				18'b000110001000011010: oled_data = 16'b1011001000101001;
				18'b000110001010011010: oled_data = 16'b1011001001001001;
				18'b000110001100011010: oled_data = 16'b1011001001001001;
				18'b000110001110011010: oled_data = 16'b1011001001001001;
				18'b000110010000011010: oled_data = 16'b1011001001001001;
				18'b000110010010011010: oled_data = 16'b1011001001001001;
				18'b000110010100011010: oled_data = 16'b1010101000101000;
				18'b000110010110011010: oled_data = 16'b1011001001001000;
				18'b000110011000011010: oled_data = 16'b1011001001001001;
				18'b000110011010011010: oled_data = 16'b1011001000101001;
				18'b000110011100011010: oled_data = 16'b1011001000101001;
				18'b000110011110011010: oled_data = 16'b1011001000101000;
				18'b000110100000011010: oled_data = 16'b1011001000101001;
				18'b000110100010011010: oled_data = 16'b1011001000101000;
				18'b000110100100011010: oled_data = 16'b1011001000101000;
				18'b000110100110011010: oled_data = 16'b1010101000101000;
				18'b000100011000011011: oled_data = 16'b0110110110111000;
				18'b000100011010011011: oled_data = 16'b0111011000111010;
				18'b000100011100011011: oled_data = 16'b0110010101011000;
				18'b000100011110011011: oled_data = 16'b0100110010010101;
				18'b000100100000011011: oled_data = 16'b0100010001110101;
				18'b000100100010011011: oled_data = 16'b0100110010110110;
				18'b000100100100011011: oled_data = 16'b0110110110111001;
				18'b000100100110011011: oled_data = 16'b0111011000111010;
				18'b000100101000011011: oled_data = 16'b1011010010110110;
				18'b000100101010011011: oled_data = 16'b1101110010010101;
				18'b000100101100011011: oled_data = 16'b1100110001110100;
				18'b000100101110011011: oled_data = 16'b1101010010010100;
				18'b000100110000011011: oled_data = 16'b1101110010110101;
				18'b000100110010011011: oled_data = 16'b1110010011010110;
				18'b000100110100011011: oled_data = 16'b1101110010010101;
				18'b000100110110011011: oled_data = 16'b1101010010010101;
				18'b000100111000011011: oled_data = 16'b1101110011010101;
				18'b000100111010011011: oled_data = 16'b1101010001110100;
				18'b000100111100011011: oled_data = 16'b1101010010010100;
				18'b000100111110011011: oled_data = 16'b1101110011010110;
				18'b000101000000011011: oled_data = 16'b1101110011010101;
				18'b000101000010011011: oled_data = 16'b1101110011010101;
				18'b000101000100011011: oled_data = 16'b1101110011010101;
				18'b000101000110011011: oled_data = 16'b1101110010110101;
				18'b000101001000011011: oled_data = 16'b1101110111010111;
				18'b000101001010011011: oled_data = 16'b1110011010011010;
				18'b000101001100011011: oled_data = 16'b1100110011010100;
				18'b000101001110011011: oled_data = 16'b1101110011010101;
				18'b000101010000011011: oled_data = 16'b1101110011010101;
				18'b000101010010011011: oled_data = 16'b1101110010110101;
				18'b000101010100011011: oled_data = 16'b1101010110010110;
				18'b000101010110011011: oled_data = 16'b1110111011111011;
				18'b000101011000011011: oled_data = 16'b1100110100010101;
				18'b000101011010011011: oled_data = 16'b1101010010010100;
				18'b000101011100011011: oled_data = 16'b1110010011010101;
				18'b000101011110011011: oled_data = 16'b1101110011010101;
				18'b000101100000011011: oled_data = 16'b1101110011010101;
				18'b000101100010011011: oled_data = 16'b1101110011010101;
				18'b000101100100011011: oled_data = 16'b1101110011010101;
				18'b000101100110011011: oled_data = 16'b1101110011010101;
				18'b000101101000011011: oled_data = 16'b1101110011010101;
				18'b000101101010011011: oled_data = 16'b1101110011010101;
				18'b000101101100011011: oled_data = 16'b1101110010110101;
				18'b000101101110011011: oled_data = 16'b1100010011010100;
				18'b000101110000011011: oled_data = 16'b0110001010101010;
				18'b000101110010011011: oled_data = 16'b0100000111000111;
				18'b000101110100011011: oled_data = 16'b1101011001111001;
				18'b000101110110011011: oled_data = 16'b1110111100011011;
				18'b000101111000011011: oled_data = 16'b1110111100011010;
				18'b000101111010011011: oled_data = 16'b1101010111110111;
				18'b000101111100011011: oled_data = 16'b1110011010111010;
				18'b000101111110011011: oled_data = 16'b1011110011010100;
				18'b000110000000011011: oled_data = 16'b1011001110110000;
				18'b000110000010011011: oled_data = 16'b1110010100010100;
				18'b000110000100011011: oled_data = 16'b1110010001110001;
				18'b000110000110011011: oled_data = 16'b1011101001101010;
				18'b000110001000011011: oled_data = 16'b1011101000101001;
				18'b000110001010011011: oled_data = 16'b1100001011101100;
				18'b000110001100011011: oled_data = 16'b1011101001101010;
				18'b000110001110011011: oled_data = 16'b1011001001001001;
				18'b000110010000011011: oled_data = 16'b1011001001001001;
				18'b000110010010011011: oled_data = 16'b1011001000101000;
				18'b000110010100011011: oled_data = 16'b1010101000101001;
				18'b000110010110011011: oled_data = 16'b1011001001001001;
				18'b000110011000011011: oled_data = 16'b1011001001001001;
				18'b000110011010011011: oled_data = 16'b1011001000001001;
				18'b000110011100011011: oled_data = 16'b1011001000101001;
				18'b000110011110011011: oled_data = 16'b1011001000101001;
				18'b000110100000011011: oled_data = 16'b1011001000101001;
				18'b000110100010011011: oled_data = 16'b1011001000101000;
				18'b000110100100011011: oled_data = 16'b1011001000101000;
				18'b000110100110011011: oled_data = 16'b1010101000101000;
				18'b000100011000011100: oled_data = 16'b0011001001101011;
				18'b000100011010011100: oled_data = 16'b0101110010010011;
				18'b000100011100011100: oled_data = 16'b0111010111111000;
				18'b000100011110011100: oled_data = 16'b0110110110111001;
				18'b000100100000011100: oled_data = 16'b0110010110111010;
				18'b000100100010011100: oled_data = 16'b0110110111111010;
				18'b000100100100011100: oled_data = 16'b0111011000111011;
				18'b000100100110011100: oled_data = 16'b0111010111111010;
				18'b000100101000011100: oled_data = 16'b1011010001110101;
				18'b000100101010011100: oled_data = 16'b1101110011010110;
				18'b000100101100011100: oled_data = 16'b1101110011010110;
				18'b000100101110011100: oled_data = 16'b1101110011110110;
				18'b000100110000011100: oled_data = 16'b1101010001110100;
				18'b000100110010011100: oled_data = 16'b1101110010110101;
				18'b000100110100011100: oled_data = 16'b1101110010110101;
				18'b000100110110011100: oled_data = 16'b1101010010010100;
				18'b000100111000011100: oled_data = 16'b1101110011010110;
				18'b000100111010011100: oled_data = 16'b1101010001110100;
				18'b000100111100011100: oled_data = 16'b1101010001110100;
				18'b000100111110011100: oled_data = 16'b1101110011010101;
				18'b000101000000011100: oled_data = 16'b1101110011010101;
				18'b000101000010011100: oled_data = 16'b1101110011010101;
				18'b000101000100011100: oled_data = 16'b1101110011010101;
				18'b000101000110011100: oled_data = 16'b1101110011010101;
				18'b000101001000011100: oled_data = 16'b1101110101110110;
				18'b000101001010011100: oled_data = 16'b1110111100011011;
				18'b000101001100011100: oled_data = 16'b1110011001111001;
				18'b000101001110011100: oled_data = 16'b1101010011010101;
				18'b000101010000011100: oled_data = 16'b1101110011010101;
				18'b000101010010011100: oled_data = 16'b1101110011010101;
				18'b000101010100011100: oled_data = 16'b1101010011010100;
				18'b000101010110011100: oled_data = 16'b1101111001111001;
				18'b000101011000011100: oled_data = 16'b1101111000111000;
				18'b000101011010011100: oled_data = 16'b1101010100010101;
				18'b000101011100011100: oled_data = 16'b1101110011010101;
				18'b000101011110011100: oled_data = 16'b1101110011010101;
				18'b000101100000011100: oled_data = 16'b1101110011010101;
				18'b000101100010011100: oled_data = 16'b1101110011010101;
				18'b000101100100011100: oled_data = 16'b1101110011010101;
				18'b000101100110011100: oled_data = 16'b1101110011010101;
				18'b000101101000011100: oled_data = 16'b1101110011010101;
				18'b000101101010011100: oled_data = 16'b1101110011010101;
				18'b000101101100011100: oled_data = 16'b1110010011010110;
				18'b000101101110011100: oled_data = 16'b1010001110110000;
				18'b000101110000011100: oled_data = 16'b0011000101000100;
				18'b000101110010011100: oled_data = 16'b1000110000010000;
				18'b000101110100011100: oled_data = 16'b1110111100011100;
				18'b000101110110011100: oled_data = 16'b1110111100011011;
				18'b000101111000011100: oled_data = 16'b1110111100111011;
				18'b000101111010011100: oled_data = 16'b1110111011011010;
				18'b000101111100011100: oled_data = 16'b1110011011011010;
				18'b000101111110011100: oled_data = 16'b1100110110110111;
				18'b000110000000011100: oled_data = 16'b1100110000110001;
				18'b000110000010011100: oled_data = 16'b1110110100010100;
				18'b000110000100011100: oled_data = 16'b1100101101101110;
				18'b000110000110011100: oled_data = 16'b1011001000101001;
				18'b000110001000011100: oled_data = 16'b1011101001101010;
				18'b000110001010011100: oled_data = 16'b1101001110001110;
				18'b000110001100011100: oled_data = 16'b1011001001101001;
				18'b000110001110011100: oled_data = 16'b1011001001001001;
				18'b000110010000011100: oled_data = 16'b1011001001001001;
				18'b000110010010011100: oled_data = 16'b1010101000001000;
				18'b000110010100011100: oled_data = 16'b1011001001001001;
				18'b000110010110011100: oled_data = 16'b1011101110001110;
				18'b000110011000011100: oled_data = 16'b1010001000101001;
				18'b000110011010011100: oled_data = 16'b1010000111000111;
				18'b000110011100011100: oled_data = 16'b1011001001001001;
				18'b000110011110011100: oled_data = 16'b1011001000101001;
				18'b000110100000011100: oled_data = 16'b1011001000101001;
				18'b000110100010011100: oled_data = 16'b1011001000101000;
				18'b000110100100011100: oled_data = 16'b1011001000101000;
				18'b000110100110011100: oled_data = 16'b1011001000101000;
				18'b000100011000011101: oled_data = 16'b0101101010101001;
				18'b000100011010011101: oled_data = 16'b1001010001001100;
				18'b000100011100011101: oled_data = 16'b1010110011010000;
				18'b000100011110011101: oled_data = 16'b1010110111010000;
				18'b000100100000011101: oled_data = 16'b1001110111110011;
				18'b000100100010011101: oled_data = 16'b1000110111110101;
				18'b000100100100011101: oled_data = 16'b1000110111110101;
				18'b000100100110011101: oled_data = 16'b1000110101110100;
				18'b000100101000011101: oled_data = 16'b1011110000010010;
				18'b000100101010011101: oled_data = 16'b1101110011010110;
				18'b000100101100011101: oled_data = 16'b1110010011110110;
				18'b000100101110011101: oled_data = 16'b1110010011010110;
				18'b000100110000011101: oled_data = 16'b1101010001010100;
				18'b000100110010011101: oled_data = 16'b1101110010110101;
				18'b000100110100011101: oled_data = 16'b1101110011010101;
				18'b000100110110011101: oled_data = 16'b1101010001110100;
				18'b000100111000011101: oled_data = 16'b1101110011010110;
				18'b000100111010011101: oled_data = 16'b1101010001110100;
				18'b000100111100011101: oled_data = 16'b1101010001110100;
				18'b000100111110011101: oled_data = 16'b1101110010110101;
				18'b000101000000011101: oled_data = 16'b1101110011010110;
				18'b000101000010011101: oled_data = 16'b1101110011010101;
				18'b000101000100011101: oled_data = 16'b1101110011010101;
				18'b000101000110011101: oled_data = 16'b1101110011010101;
				18'b000101001000011101: oled_data = 16'b1101010100110110;
				18'b000101001010011101: oled_data = 16'b1110111100011011;
				18'b000101001100011101: oled_data = 16'b1110111100011011;
				18'b000101001110011101: oled_data = 16'b1101111001111001;
				18'b000101010000011101: oled_data = 16'b1101010011010101;
				18'b000101010010011101: oled_data = 16'b1101110011010101;
				18'b000101010100011101: oled_data = 16'b1101110011010101;
				18'b000101010110011101: oled_data = 16'b1100110100010101;
				18'b000101011000011101: oled_data = 16'b1110011011111010;
				18'b000101011010011101: oled_data = 16'b1110011011011010;
				18'b000101011100011101: oled_data = 16'b1101010100110101;
				18'b000101011110011101: oled_data = 16'b1101110011010101;
				18'b000101100000011101: oled_data = 16'b1101110011010101;
				18'b000101100010011101: oled_data = 16'b1101110011010101;
				18'b000101100100011101: oled_data = 16'b1101110011010101;
				18'b000101100110011101: oled_data = 16'b1101110011010101;
				18'b000101101000011101: oled_data = 16'b1101110011010101;
				18'b000101101010011101: oled_data = 16'b1101110011010101;
				18'b000101101100011101: oled_data = 16'b1110010011110110;
				18'b000101101110011101: oled_data = 16'b0111101010001011;
				18'b000101110000011101: oled_data = 16'b0100000111000110;
				18'b000101110010011101: oled_data = 16'b1101011001111001;
				18'b000101110100011101: oled_data = 16'b1111011100111100;
				18'b000101110110011101: oled_data = 16'b1101111010011001;
				18'b000101111000011101: oled_data = 16'b1011010100110100;
				18'b000101111010011101: oled_data = 16'b0111101101001101;
				18'b000101111100011101: oled_data = 16'b1010110100010011;
				18'b000101111110011101: oled_data = 16'b1100110111010110;
				18'b000110000000011101: oled_data = 16'b1110010011010100;
				18'b000110000010011101: oled_data = 16'b1110010011010011;
				18'b000110000100011101: oled_data = 16'b1011101010001010;
				18'b000110000110011101: oled_data = 16'b1011101000101001;
				18'b000110001000011101: oled_data = 16'b1100001011001011;
				18'b000110001010011101: oled_data = 16'b1100001100101100;
				18'b000110001100011101: oled_data = 16'b1011001001001001;
				18'b000110001110011101: oled_data = 16'b1011001001001001;
				18'b000110010000011101: oled_data = 16'b1010101000101000;
				18'b000110010010011101: oled_data = 16'b1011001000101001;
				18'b000110010100011101: oled_data = 16'b1011001010001011;
				18'b000110010110011101: oled_data = 16'b1011111000111000;
				18'b000110011000011101: oled_data = 16'b1010001101001101;
				18'b000110011010011101: oled_data = 16'b1010100111101000;
				18'b000110011100011101: oled_data = 16'b1011001001001001;
				18'b000110011110011101: oled_data = 16'b1011001000101001;
				18'b000110100000011101: oled_data = 16'b1011001000101001;
				18'b000110100010011101: oled_data = 16'b1011001000101000;
				18'b000110100100011101: oled_data = 16'b1011001000101000;
				18'b000110100110011101: oled_data = 16'b1011001000101000;
				18'b000100011000011110: oled_data = 16'b1100110011001111;
				18'b000100011010011110: oled_data = 16'b1100110011110001;
				18'b000100011100011110: oled_data = 16'b1101011000101110;
				18'b000100011110011110: oled_data = 16'b1110011011010001;
				18'b000100100000011110: oled_data = 16'b1110011011110010;
				18'b000100100010011110: oled_data = 16'b1101011000101101;
				18'b000100100100011110: oled_data = 16'b1100110111001010;
				18'b000100100110011110: oled_data = 16'b1101010111101100;
				18'b000100101000011110: oled_data = 16'b1011110000110000;
				18'b000100101010011110: oled_data = 16'b1101010001110101;
				18'b000100101100011110: oled_data = 16'b1101110011010101;
				18'b000100101110011110: oled_data = 16'b1110010011010110;
				18'b000100110000011110: oled_data = 16'b1100110000110011;
				18'b000100110010011110: oled_data = 16'b1101010001110100;
				18'b000100110100011110: oled_data = 16'b1110010011010110;
				18'b000100110110011110: oled_data = 16'b1101010001110100;
				18'b000100111000011110: oled_data = 16'b1101110011010101;
				18'b000100111010011110: oled_data = 16'b1101010010010100;
				18'b000100111100011110: oled_data = 16'b1101010010010101;
				18'b000100111110011110: oled_data = 16'b1101010010010100;
				18'b000101000000011110: oled_data = 16'b1101110011010110;
				18'b000101000010011110: oled_data = 16'b1101110011010101;
				18'b000101000100011110: oled_data = 16'b1101110011010101;
				18'b000101000110011110: oled_data = 16'b1110010011010110;
				18'b000101001000011110: oled_data = 16'b1101010100110101;
				18'b000101001010011110: oled_data = 16'b1110011100011010;
				18'b000101001100011110: oled_data = 16'b1110011100011010;
				18'b000101001110011110: oled_data = 16'b1110111100111011;
				18'b000101010000011110: oled_data = 16'b1101111000011001;
				18'b000101010010011110: oled_data = 16'b1100110010010100;
				18'b000101010100011110: oled_data = 16'b1101010010010100;
				18'b000101010110011110: oled_data = 16'b1101010011010100;
				18'b000101011000011110: oled_data = 16'b1101111001111000;
				18'b000101011010011110: oled_data = 16'b1110111100111011;
				18'b000101011100011110: oled_data = 16'b1101111011011010;
				18'b000101011110011110: oled_data = 16'b1101010100110110;
				18'b000101100000011110: oled_data = 16'b1101110010110101;
				18'b000101100010011110: oled_data = 16'b1101110011010101;
				18'b000101100100011110: oled_data = 16'b1101110011010101;
				18'b000101100110011110: oled_data = 16'b1101110011010101;
				18'b000101101000011110: oled_data = 16'b1101110011010101;
				18'b000101101010011110: oled_data = 16'b1101110011010110;
				18'b000101101100011110: oled_data = 16'b1101010001110100;
				18'b000101101110011110: oled_data = 16'b0101000110000111;
				18'b000101110000011110: oled_data = 16'b0111001101001100;
				18'b000101110010011110: oled_data = 16'b1011010100110100;
				18'b000101110100011110: oled_data = 16'b0111001100101100;
				18'b000101110110011110: oled_data = 16'b0100000110100110;
				18'b000101111000011110: oled_data = 16'b0100000110100110;
				18'b000101111010011110: oled_data = 16'b1000001111101111;
				18'b000101111100011110: oled_data = 16'b1100111000110111;
				18'b000101111110011110: oled_data = 16'b1100110101110101;
				18'b000110000000011110: oled_data = 16'b1110110011110100;
				18'b000110000010011110: oled_data = 16'b1101001111110000;
				18'b000110000100011110: oled_data = 16'b1010101000101000;
				18'b000110000110011110: oled_data = 16'b1011101000101001;
				18'b000110001000011110: oled_data = 16'b1100101100001100;
				18'b000110001010011110: oled_data = 16'b1011101010101010;
				18'b000110001100011110: oled_data = 16'b1011001001001001;
				18'b000110001110011110: oled_data = 16'b1011001001001001;
				18'b000110010000011110: oled_data = 16'b1010101000101000;
				18'b000110010010011110: oled_data = 16'b1011101001001001;
				18'b000110010100011110: oled_data = 16'b1011101110101111;
				18'b000110010110011110: oled_data = 16'b1011111100011100;
				18'b000110011000011110: oled_data = 16'b1011010101110110;
				18'b000110011010011110: oled_data = 16'b1011001010001010;
				18'b000110011100011110: oled_data = 16'b1011101010101010;
				18'b000110011110011110: oled_data = 16'b1011001000101000;
				18'b000110100000011110: oled_data = 16'b1011001000101001;
				18'b000110100010011110: oled_data = 16'b1011001000101001;
				18'b000110100100011110: oled_data = 16'b1011001000001000;
				18'b000110100110011110: oled_data = 16'b1010101000001000;
				18'b000100011000011111: oled_data = 16'b1101010011110010;
				18'b000100011010011111: oled_data = 16'b1101111000010001;
				18'b000100011100011111: oled_data = 16'b1110111100010101;
				18'b000100011110011111: oled_data = 16'b1110011011010101;
				18'b000100100000011111: oled_data = 16'b1110011011010100;
				18'b000100100010011111: oled_data = 16'b1101011000010000;
				18'b000100100100011111: oled_data = 16'b1010110011001000;
				18'b000100100110011111: oled_data = 16'b1100110111101011;
				18'b000100101000011111: oled_data = 16'b1100110011110000;
				18'b000100101010011111: oled_data = 16'b1101110010110110;
				18'b000100101100011111: oled_data = 16'b1101010001110100;
				18'b000100101110011111: oled_data = 16'b1101110011010101;
				18'b000100110000011111: oled_data = 16'b1100110000110011;
				18'b000100110010011111: oled_data = 16'b1100110000110011;
				18'b000100110100011111: oled_data = 16'b1110010011110110;
				18'b000100110110011111: oled_data = 16'b1101010010010100;
				18'b000100111000011111: oled_data = 16'b1101110010110101;
				18'b000100111010011111: oled_data = 16'b1101110010010101;
				18'b000100111100011111: oled_data = 16'b1101110010010101;
				18'b000100111110011111: oled_data = 16'b1101010001110100;
				18'b000101000000011111: oled_data = 16'b1101110011010101;
				18'b000101000010011111: oled_data = 16'b1101110011010101;
				18'b000101000100011111: oled_data = 16'b1101110011010101;
				18'b000101000110011111: oled_data = 16'b1110010011010110;
				18'b000101001000011111: oled_data = 16'b1100110011110101;
				18'b000101001010011111: oled_data = 16'b1110011011111010;
				18'b000101001100011111: oled_data = 16'b1110111100011010;
				18'b000101001110011111: oled_data = 16'b1110111100011010;
				18'b000101010000011111: oled_data = 16'b1101111010111001;
				18'b000101010010011111: oled_data = 16'b1100110110110110;
				18'b000101010100011111: oled_data = 16'b1101010011010101;
				18'b000101010110011111: oled_data = 16'b1101110011110101;
				18'b000101011000011111: oled_data = 16'b1101010101010110;
				18'b000101011010011111: oled_data = 16'b1110111011111011;
				18'b000101011100011111: oled_data = 16'b1110111100011011;
				18'b000101011110011111: oled_data = 16'b1110011010111010;
				18'b000101100000011111: oled_data = 16'b1101010101010110;
				18'b000101100010011111: oled_data = 16'b1101110010110101;
				18'b000101100100011111: oled_data = 16'b1101110011010101;
				18'b000101100110011111: oled_data = 16'b1101110011010101;
				18'b000101101000011111: oled_data = 16'b1101110011010101;
				18'b000101101010011111: oled_data = 16'b1110010011110110;
				18'b000101101100011111: oled_data = 16'b1011001110010000;
				18'b000101101110011111: oled_data = 16'b0100100101100110;
				18'b000101110000011111: oled_data = 16'b0011100101000101;
				18'b000101110010011111: oled_data = 16'b0011000100100100;
				18'b000101110100011111: oled_data = 16'b0100100111100111;
				18'b000101110110011111: oled_data = 16'b1000001111001111;
				18'b000101111000011111: oled_data = 16'b1100111000111000;
				18'b000101111010011111: oled_data = 16'b1110111100111100;
				18'b000101111100011111: oled_data = 16'b1101011001111000;
				18'b000101111110011111: oled_data = 16'b1101010100110100;
				18'b000110000000011111: oled_data = 16'b1110110011110100;
				18'b000110000010011111: oled_data = 16'b1100001100001101;
				18'b000110000100011111: oled_data = 16'b1011001000101000;
				18'b000110000110011111: oled_data = 16'b1011101001001001;
				18'b000110001000011111: oled_data = 16'b1011101010001010;
				18'b000110001010011111: oled_data = 16'b1011101001001001;
				18'b000110001100011111: oled_data = 16'b1011001001001001;
				18'b000110001110011111: oled_data = 16'b1010101000001000;
				18'b000110010000011111: oled_data = 16'b1011001000101001;
				18'b000110010010011111: oled_data = 16'b1011001000001001;
				18'b000110010100011111: oled_data = 16'b1011110101010110;
				18'b000110010110011111: oled_data = 16'b1011111100011100;
				18'b000110011000011111: oled_data = 16'b1011111010111011;
				18'b000110011010011111: oled_data = 16'b1101010001010010;
				18'b000110011100011111: oled_data = 16'b1011101010001010;
				18'b000110011110011111: oled_data = 16'b1011001000101001;
				18'b000110100000011111: oled_data = 16'b1011001000101001;
				18'b000110100010011111: oled_data = 16'b1011001000101000;
				18'b000110100100011111: oled_data = 16'b1011001000001000;
				18'b000110100110011111: oled_data = 16'b1010101000001000;
				18'b000100011000100000: oled_data = 16'b1100110110001101;
				18'b000100011010100000: oled_data = 16'b1100010110101100;
				18'b000100011100100000: oled_data = 16'b1011110101101100;
				18'b000100011110100000: oled_data = 16'b1010110011101001;
				18'b000100100000100000: oled_data = 16'b1010110011001000;
				18'b000100100010100000: oled_data = 16'b1100110110101101;
				18'b000100100100100000: oled_data = 16'b1010110011001000;
				18'b000100100110100000: oled_data = 16'b1011010100101001;
				18'b000100101000100000: oled_data = 16'b1101010101101111;
				18'b000100101010100000: oled_data = 16'b1101110011010101;
				18'b000100101100100000: oled_data = 16'b1101110011010110;
				18'b000100101110100000: oled_data = 16'b1101110011010101;
				18'b000100110000100000: oled_data = 16'b1100110000110011;
				18'b000100110010100000: oled_data = 16'b1100001111110010;
				18'b000100110100100000: oled_data = 16'b1110010011110110;
				18'b000100110110100000: oled_data = 16'b1101110010110101;
				18'b000100111000100000: oled_data = 16'b1101010010010101;
				18'b000100111010100000: oled_data = 16'b1101110010110101;
				18'b000100111100100000: oled_data = 16'b1101010010010101;
				18'b000100111110100000: oled_data = 16'b1101010010010100;
				18'b000101000000100000: oled_data = 16'b1101110010110101;
				18'b000101000010100000: oled_data = 16'b1101110011010110;
				18'b000101000100100000: oled_data = 16'b1101110011010101;
				18'b000101000110100000: oled_data = 16'b1110010011010110;
				18'b000101001000100000: oled_data = 16'b1100110011110101;
				18'b000101001010100000: oled_data = 16'b1110011011011010;
				18'b000101001100100000: oled_data = 16'b1101111010111001;
				18'b000101001110100000: oled_data = 16'b1101111010111001;
				18'b000101010000100000: oled_data = 16'b1110011011111010;
				18'b000101010010100000: oled_data = 16'b1110111100111011;
				18'b000101010100100000: oled_data = 16'b1110011000111000;
				18'b000101010110100000: oled_data = 16'b1101010100010101;
				18'b000101011000100000: oled_data = 16'b1101110011010101;
				18'b000101011010100000: oled_data = 16'b1101110111111001;
				18'b000101011100100000: oled_data = 16'b1110111100011011;
				18'b000101011110100000: oled_data = 16'b1110111100011010;
				18'b000101100000100000: oled_data = 16'b1110011011011010;
				18'b000101100010100000: oled_data = 16'b1101110110010111;
				18'b000101100100100000: oled_data = 16'b1101110010110101;
				18'b000101100110100000: oled_data = 16'b1110010011010101;
				18'b000101101000100000: oled_data = 16'b1101110011010110;
				18'b000101101010100000: oled_data = 16'b1101110011010110;
				18'b000101101100100000: oled_data = 16'b1000101010101100;
				18'b000101101110100000: oled_data = 16'b0101000111101000;
				18'b000101110000100000: oled_data = 16'b0111101110001110;
				18'b000101110010100000: oled_data = 16'b1011010101010101;
				18'b000101110100100000: oled_data = 16'b1101111010111010;
				18'b000101110110100000: oled_data = 16'b1110111100111100;
				18'b000101111000100000: oled_data = 16'b1110111100011011;
				18'b000101111010100000: oled_data = 16'b1101111011011010;
				18'b000101111100100000: oled_data = 16'b1101011000110111;
				18'b000101111110100000: oled_data = 16'b1101110100010100;
				18'b000110000000100000: oled_data = 16'b1110010011010011;
				18'b000110000010100000: oled_data = 16'b1011001010001010;
				18'b000110000100100000: oled_data = 16'b1011001000101001;
				18'b000110000110100000: oled_data = 16'b1011101001001001;
				18'b000110001000100000: oled_data = 16'b1011101000101001;
				18'b000110001010100000: oled_data = 16'b1011001001001001;
				18'b000110001100100000: oled_data = 16'b1011001001001001;
				18'b000110001110100000: oled_data = 16'b1011001000001000;
				18'b000110010000100000: oled_data = 16'b1011001000001001;
				18'b000110010010100000: oled_data = 16'b1010101011001100;
				18'b000110010100100000: oled_data = 16'b1011111010111010;
				18'b000110010110100000: oled_data = 16'b1011111011111011;
				18'b000110011000100000: oled_data = 16'b1011111100011100;
				18'b000110011010100000: oled_data = 16'b1011110100110101;
				18'b000110011100100000: oled_data = 16'b1011001000001001;
				18'b000110011110100000: oled_data = 16'b1011001000101001;
				18'b000110100000100000: oled_data = 16'b1011001000101000;
				18'b000110100010100000: oled_data = 16'b1011001000101000;
				18'b000110100100100000: oled_data = 16'b1011001000001000;
				18'b000110100110100000: oled_data = 16'b1010101000001000;
				18'b000100011000100001: oled_data = 16'b1100110111001100;
				18'b000100011010100001: oled_data = 16'b1010110011001000;
				18'b000100011100100001: oled_data = 16'b1010110010100111;
				18'b000100011110100001: oled_data = 16'b1010110010100111;
				18'b000100100000100001: oled_data = 16'b1010110010100111;
				18'b000100100010100001: oled_data = 16'b1011110101001011;
				18'b000100100100100001: oled_data = 16'b1010110011001000;
				18'b000100100110100001: oled_data = 16'b1010110011101000;
				18'b000100101000100001: oled_data = 16'b1101010110001101;
				18'b000100101010100001: oled_data = 16'b1101110010110101;
				18'b000100101100100001: oled_data = 16'b1101010010010101;
				18'b000100101110100001: oled_data = 16'b1101110011010101;
				18'b000100110000100001: oled_data = 16'b1100110000110011;
				18'b000100110010100001: oled_data = 16'b1011101110110001;
				18'b000100110100100001: oled_data = 16'b1101110011010101;
				18'b000100110110100001: oled_data = 16'b1101110011010101;
				18'b000100111000100001: oled_data = 16'b1101010001110100;
				18'b000100111010100001: oled_data = 16'b1101110010110101;
				18'b000100111100100001: oled_data = 16'b1101010001110100;
				18'b000100111110100001: oled_data = 16'b1101110010110101;
				18'b000101000000100001: oled_data = 16'b1101010001110100;
				18'b000101000010100001: oled_data = 16'b1101110011010110;
				18'b000101000100100001: oled_data = 16'b1101110011010101;
				18'b000101000110100001: oled_data = 16'b1110010011010110;
				18'b000101001000100001: oled_data = 16'b1100110011110101;
				18'b000101001010100001: oled_data = 16'b1101011001011000;
				18'b000101001100100001: oled_data = 16'b1101111011011001;
				18'b000101001110100001: oled_data = 16'b1110111100011010;
				18'b000101010000100001: oled_data = 16'b1110111100011010;
				18'b000101010010100001: oled_data = 16'b1110111100011010;
				18'b000101010100100001: oled_data = 16'b1110111100111011;
				18'b000101010110100001: oled_data = 16'b1110011010111001;
				18'b000101011000100001: oled_data = 16'b1101010101010110;
				18'b000101011010100001: oled_data = 16'b1101010011110101;
				18'b000101011100100001: oled_data = 16'b1110011010111010;
				18'b000101011110100001: oled_data = 16'b1110111100011010;
				18'b000101100000100001: oled_data = 16'b1110111100011010;
				18'b000101100010100001: oled_data = 16'b1110111011111011;
				18'b000101100100100001: oled_data = 16'b1110011000011000;
				18'b000101100110100001: oled_data = 16'b1101010011110101;
				18'b000101101000100001: oled_data = 16'b1101010011010101;
				18'b000101101010100001: oled_data = 16'b1101110011010101;
				18'b000101101100100001: oled_data = 16'b1100010000110011;
				18'b000101101110100001: oled_data = 16'b1100110110010110;
				18'b000101110000100001: oled_data = 16'b1111011100111100;
				18'b000101110010100001: oled_data = 16'b1110111100111011;
				18'b000101110100100001: oled_data = 16'b1110111100011011;
				18'b000101110110100001: oled_data = 16'b1110111100011011;
				18'b000101111000100001: oled_data = 16'b1110011011111010;
				18'b000101111010100001: oled_data = 16'b1101011010011000;
				18'b000101111100100001: oled_data = 16'b1101111000010111;
				18'b000101111110100001: oled_data = 16'b1110010100010100;
				18'b000110000000100001: oled_data = 16'b1101110001110001;
				18'b000110000010100001: oled_data = 16'b1010101000101001;
				18'b000110000100100001: oled_data = 16'b1011001001001001;
				18'b000110000110100001: oled_data = 16'b1011001001001001;
				18'b000110001000100001: oled_data = 16'b1011001001001001;
				18'b000110001010100001: oled_data = 16'b1011001001001001;
				18'b000110001100100001: oled_data = 16'b1010101000101000;
				18'b000110001110100001: oled_data = 16'b1011001001001001;
				18'b000110010000100001: oled_data = 16'b1010100111001000;
				18'b000110010010100001: oled_data = 16'b1011010010110010;
				18'b000110010100100001: oled_data = 16'b1100011100011100;
				18'b000110010110100001: oled_data = 16'b1011111011111011;
				18'b000110011000100001: oled_data = 16'b1011111011111100;
				18'b000110011010100001: oled_data = 16'b1011111010011010;
				18'b000110011100100001: oled_data = 16'b1011001011101100;
				18'b000110011110100001: oled_data = 16'b1011001000101001;
				18'b000110100000100001: oled_data = 16'b1011001000101001;
				18'b000110100010100001: oled_data = 16'b1011001000101000;
				18'b000110100100100001: oled_data = 16'b1011001000001000;
				18'b000110100110100001: oled_data = 16'b1010101000001000;
				18'b000100011000100010: oled_data = 16'b1100010110101011;
				18'b000100011010100010: oled_data = 16'b1011010011101000;
				18'b000100011100100010: oled_data = 16'b1010110010100111;
				18'b000100011110100010: oled_data = 16'b1010110010100111;
				18'b000100100000100010: oled_data = 16'b1010110010100111;
				18'b000100100010100010: oled_data = 16'b1011110100101011;
				18'b000100100100100010: oled_data = 16'b1010110011101000;
				18'b000100100110100010: oled_data = 16'b1010110011001000;
				18'b000100101000100010: oled_data = 16'b1101010110101100;
				18'b000100101010100010: oled_data = 16'b1101110011010101;
				18'b000100101100100010: oled_data = 16'b1100110000010011;
				18'b000100101110100010: oled_data = 16'b1011101111010001;
				18'b000100110000100010: oled_data = 16'b1011101111010001;
				18'b000100110010100010: oled_data = 16'b1011001110010001;
				18'b000100110100100010: oled_data = 16'b1101110010110101;
				18'b000100110110100010: oled_data = 16'b1110010011010110;
				18'b000100111000100010: oled_data = 16'b1101010010010100;
				18'b000100111010100010: oled_data = 16'b1101010010010101;
				18'b000100111100100010: oled_data = 16'b1101010001110100;
				18'b000100111110100010: oled_data = 16'b1101110011010101;
				18'b000101000000100010: oled_data = 16'b1101010001110100;
				18'b000101000010100010: oled_data = 16'b1101110010110101;
				18'b000101000100100010: oled_data = 16'b1101110011010110;
				18'b000101000110100010: oled_data = 16'b1101110011010101;
				18'b000101001000100010: oled_data = 16'b1101010100110110;
				18'b000101001010100010: oled_data = 16'b1110011100011010;
				18'b000101001100100010: oled_data = 16'b1110111100011010;
				18'b000101001110100010: oled_data = 16'b1110111100011010;
				18'b000101010000100010: oled_data = 16'b1110111100011010;
				18'b000101010010100010: oled_data = 16'b1110111100011010;
				18'b000101010100100010: oled_data = 16'b1110111100011010;
				18'b000101010110100010: oled_data = 16'b1110111100111010;
				18'b000101011000100010: oled_data = 16'b1110111011111010;
				18'b000101011010100010: oled_data = 16'b1101010111110111;
				18'b000101011100100010: oled_data = 16'b1100010110110110;
				18'b000101011110100010: oled_data = 16'b1110111011111010;
				18'b000101100000100010: oled_data = 16'b1110111100011010;
				18'b000101100010100010: oled_data = 16'b1110111100011010;
				18'b000101100100100010: oled_data = 16'b1110111100011010;
				18'b000101100110100010: oled_data = 16'b1110011011011010;
				18'b000101101000100010: oled_data = 16'b1101010110110110;
				18'b000101101010100010: oled_data = 16'b1101010011110100;
				18'b000101101100100010: oled_data = 16'b1101110010010100;
				18'b000101101110100010: oled_data = 16'b1101111000011000;
				18'b000101110000100010: oled_data = 16'b1110111100011010;
				18'b000101110010100010: oled_data = 16'b1110111100011010;
				18'b000101110100100010: oled_data = 16'b1110111100011010;
				18'b000101110110100010: oled_data = 16'b1110111100011010;
				18'b000101111000100010: oled_data = 16'b1101111010111001;
				18'b000101111010100010: oled_data = 16'b1101111011111001;
				18'b000101111100100010: oled_data = 16'b1101110110110110;
				18'b000101111110100010: oled_data = 16'b1110010100010100;
				18'b000110000000100010: oled_data = 16'b1100101110101111;
				18'b000110000010100010: oled_data = 16'b1010101000101000;
				18'b000110000100100010: oled_data = 16'b1011001001001001;
				18'b000110000110100010: oled_data = 16'b1011001001001001;
				18'b000110001000100010: oled_data = 16'b1011001001001001;
				18'b000110001010100010: oled_data = 16'b1011001001001001;
				18'b000110001100100010: oled_data = 16'b1010101000101000;
				18'b000110001110100010: oled_data = 16'b1011001000101001;
				18'b000110010000100010: oled_data = 16'b1001101000101001;
				18'b000110010010100010: oled_data = 16'b1011111001111001;
				18'b000110010100100010: oled_data = 16'b1011111011111100;
				18'b000110010110100010: oled_data = 16'b1011111011111011;
				18'b000110011000100010: oled_data = 16'b1011111011111011;
				18'b000110011010100010: oled_data = 16'b1100011100011100;
				18'b000110011100100010: oled_data = 16'b1011110001110010;
				18'b000110011110100010: oled_data = 16'b1011001000001000;
				18'b000110100000100010: oled_data = 16'b1011001000101001;
				18'b000110100010100010: oled_data = 16'b1011001000101000;
				18'b000110100100100010: oled_data = 16'b1011001000001000;
				18'b000110100110100010: oled_data = 16'b1010101000001000;
				18'b000100011000100011: oled_data = 16'b1011010101001011;
				18'b000100011010100011: oled_data = 16'b1011010011101000;
				18'b000100011100100011: oled_data = 16'b1010110010100111;
				18'b000100011110100011: oled_data = 16'b1010110010100111;
				18'b000100100000100011: oled_data = 16'b1010110010100111;
				18'b000100100010100011: oled_data = 16'b1011010011101001;
				18'b000100100100100011: oled_data = 16'b1010110011001000;
				18'b000100100110100011: oled_data = 16'b1010110011000111;
				18'b000100101000100011: oled_data = 16'b1101010111001100;
				18'b000100101010100011: oled_data = 16'b1101110011110101;
				18'b000100101100100011: oled_data = 16'b1101110010110101;
				18'b000100101110100011: oled_data = 16'b1100001111010010;
				18'b000100110000100011: oled_data = 16'b1011001110010000;
				18'b000100110010100011: oled_data = 16'b1011001101110000;
				18'b000100110100100011: oled_data = 16'b1101110010110101;
				18'b000100110110100011: oled_data = 16'b1101110011010110;
				18'b000100111000100011: oled_data = 16'b1101110010110101;
				18'b000100111010100011: oled_data = 16'b1101010001110100;
				18'b000100111100100011: oled_data = 16'b1101010010010100;
				18'b000100111110100011: oled_data = 16'b1101110011010101;
				18'b000101000000100011: oled_data = 16'b1101110010110101;
				18'b000101000010100011: oled_data = 16'b1101010001110100;
				18'b000101000100100011: oled_data = 16'b1101110011010101;
				18'b000101000110100011: oled_data = 16'b1101110011010101;
				18'b000101001000100011: oled_data = 16'b1101010101110110;
				18'b000101001010100011: oled_data = 16'b1110111100111011;
				18'b000101001100100011: oled_data = 16'b1110111100011010;
				18'b000101001110100011: oled_data = 16'b1110111100111011;
				18'b000101010000100011: oled_data = 16'b1110111100111011;
				18'b000101010010100011: oled_data = 16'b1111011100111011;
				18'b000101010100100011: oled_data = 16'b1111011101011011;
				18'b000101010110100011: oled_data = 16'b1111011101011011;
				18'b000101011000100011: oled_data = 16'b1111011100111011;
				18'b000101011010100011: oled_data = 16'b1110111100011011;
				18'b000101011100100011: oled_data = 16'b1101011001111000;
				18'b000101011110100011: oled_data = 16'b1101011001011000;
				18'b000101100000100011: oled_data = 16'b1101111010111001;
				18'b000101100010100011: oled_data = 16'b1110111100011010;
				18'b000101100100100011: oled_data = 16'b1110111100011010;
				18'b000101100110100011: oled_data = 16'b1110111100011011;
				18'b000101101000100011: oled_data = 16'b1110111100111011;
				18'b000101101010100011: oled_data = 16'b1110011010111010;
				18'b000101101100100011: oled_data = 16'b1101010110110111;
				18'b000101101110100011: oled_data = 16'b1110011001111001;
				18'b000101110000100011: oled_data = 16'b1110111100011010;
				18'b000101110010100011: oled_data = 16'b1110111100011010;
				18'b000101110100100011: oled_data = 16'b1110111100011010;
				18'b000101110110100011: oled_data = 16'b1110011011111010;
				18'b000101111000100011: oled_data = 16'b1101111010011000;
				18'b000101111010100011: oled_data = 16'b1110011100011010;
				18'b000101111100100011: oled_data = 16'b1101010101110101;
				18'b000101111110100011: oled_data = 16'b1110110011110100;
				18'b000110000000100011: oled_data = 16'b1011101100101100;
				18'b000110000010100011: oled_data = 16'b1010101000101000;
				18'b000110000100100011: oled_data = 16'b1011001001001001;
				18'b000110000110100011: oled_data = 16'b1011001001001001;
				18'b000110001000100011: oled_data = 16'b1011101001001001;
				18'b000110001010100011: oled_data = 16'b1011001000101001;
				18'b000110001100100011: oled_data = 16'b1010101000101001;
				18'b000110001110100011: oled_data = 16'b1010000111001000;
				18'b000110010000100011: oled_data = 16'b1010001110001111;
				18'b000110010010100011: oled_data = 16'b1011111100011011;
				18'b000110010100100011: oled_data = 16'b1011111011111011;
				18'b000110010110100011: oled_data = 16'b1011111011111011;
				18'b000110011000100011: oled_data = 16'b1011111011111011;
				18'b000110011010100011: oled_data = 16'b1100111100111100;
				18'b000110011100100011: oled_data = 16'b1011111000010111;
				18'b000110011110100011: oled_data = 16'b1011001001101001;
				18'b000110100000100011: oled_data = 16'b1011001000101001;
				18'b000110100010100011: oled_data = 16'b1011001000101001;
				18'b000110100100100011: oled_data = 16'b1011001000001000;
				18'b000110100110100011: oled_data = 16'b1010101000001000;
				18'b000100011000100100: oled_data = 16'b1001110010101010;
				18'b000100011010100100: oled_data = 16'b1100010101001001;
				18'b000100011100100100: oled_data = 16'b1010110010000111;
				18'b000100011110100100: oled_data = 16'b1010110010100111;
				18'b000100100000100100: oled_data = 16'b1010110010100111;
				18'b000100100010100100: oled_data = 16'b1010110010100111;
				18'b000100100100100100: oled_data = 16'b1010110010000111;
				18'b000100100110100100: oled_data = 16'b1011010100001000;
				18'b000100101000100100: oled_data = 16'b1101011000001100;
				18'b000100101010100100: oled_data = 16'b1101110011110100;
				18'b000100101100100100: oled_data = 16'b1110010011010110;
				18'b000100101110100100: oled_data = 16'b1101010010110101;
				18'b000100110000100100: oled_data = 16'b1011001111010001;
				18'b000100110010100100: oled_data = 16'b1010101101010000;
				18'b000100110100100100: oled_data = 16'b1101010010010101;
				18'b000100110110100100: oled_data = 16'b1101110011010110;
				18'b000100111000100100: oled_data = 16'b1101110011010110;
				18'b000100111010100100: oled_data = 16'b1101010010010100;
				18'b000100111100100100: oled_data = 16'b1100110001010011;
				18'b000100111110100100: oled_data = 16'b1101110011010101;
				18'b000101000000100100: oled_data = 16'b1101110011010101;
				18'b000101000010100100: oled_data = 16'b1101110010010101;
				18'b000101000100100100: oled_data = 16'b1101010010010100;
				18'b000101000110100100: oled_data = 16'b1110010011110110;
				18'b000101001000100100: oled_data = 16'b1101110110110111;
				18'b000101001010100100: oled_data = 16'b1110111100011011;
				18'b000101001100100100: oled_data = 16'b1110011011011001;
				18'b000101001110100100: oled_data = 16'b1101011001111000;
				18'b000101010000100100: oled_data = 16'b1100111000010111;
				18'b000101010010100100: oled_data = 16'b1011010101010100;
				18'b000101010100100100: oled_data = 16'b1001110010010001;
				18'b000101010110100100: oled_data = 16'b1000110000001111;
				18'b000101011000100100: oled_data = 16'b0111001101001100;
				18'b000101011010100100: oled_data = 16'b0110001011001010;
				18'b000101011100100100: oled_data = 16'b0101001001101001;
				18'b000101011110100100: oled_data = 16'b0011100110100110;
				18'b000101100000100100: oled_data = 16'b1001010001110000;
				18'b000101100010100100: oled_data = 16'b1110111101011011;
				18'b000101100100100100: oled_data = 16'b1110111100011010;
				18'b000101100110100100: oled_data = 16'b1110111100011010;
				18'b000101101000100100: oled_data = 16'b1110111100011010;
				18'b000101101010100100: oled_data = 16'b1110011100111011;
				18'b000101101100100100: oled_data = 16'b1110111100111011;
				18'b000101101110100100: oled_data = 16'b1110111100011011;
				18'b000101110000100100: oled_data = 16'b1110111100011010;
				18'b000101110010100100: oled_data = 16'b1110111100011010;
				18'b000101110100100100: oled_data = 16'b1110111100011010;
				18'b000101110110100100: oled_data = 16'b1101111010011000;
				18'b000101111000100100: oled_data = 16'b1110011011111010;
				18'b000101111010100100: oled_data = 16'b1110011011111010;
				18'b000101111100100100: oled_data = 16'b1101010101010100;
				18'b000101111110100100: oled_data = 16'b1110110011110011;
				18'b000110000000100100: oled_data = 16'b1011101010101011;
				18'b000110000010100100: oled_data = 16'b1011001000101001;
				18'b000110000100100100: oled_data = 16'b1011001001001001;
				18'b000110000110100100: oled_data = 16'b1011001001001001;
				18'b000110001000100100: oled_data = 16'b1011101000101001;
				18'b000110001010100100: oled_data = 16'b1010101000001000;
				18'b000110001100100100: oled_data = 16'b1010101000101001;
				18'b000110001110100100: oled_data = 16'b1001100110000111;
				18'b000110010000100100: oled_data = 16'b1011010100110101;
				18'b000110010010100100: oled_data = 16'b1011111100011100;
				18'b000110010100100100: oled_data = 16'b1011111011111011;
				18'b000110010110100100: oled_data = 16'b1011111011111011;
				18'b000110011000100100: oled_data = 16'b1011111011111011;
				18'b000110011010100100: oled_data = 16'b1100111100011100;
				18'b000110011100100100: oled_data = 16'b1011111011111011;
				18'b000110011110100100: oled_data = 16'b1011001100101101;
				18'b000110100000100100: oled_data = 16'b1011001000001000;
				18'b000110100010100100: oled_data = 16'b1011001000101001;
				18'b000110100100100100: oled_data = 16'b1010101000101000;
				18'b000110100110100100: oled_data = 16'b1010101000101000;
				18'b000100011000100101: oled_data = 16'b1000001111001000;
				18'b000100011010100101: oled_data = 16'b1101011000101011;
				18'b000100011100100101: oled_data = 16'b1011010011101000;
				18'b000100011110100101: oled_data = 16'b1010110010100111;
				18'b000100100000100101: oled_data = 16'b1010110010100111;
				18'b000100100010100101: oled_data = 16'b1010110010000111;
				18'b000100100100100101: oled_data = 16'b1010110010100111;
				18'b000100100110100101: oled_data = 16'b1100110111001010;
				18'b000100101000100101: oled_data = 16'b1101111000001100;
				18'b000100101010100101: oled_data = 16'b1101110011010100;
				18'b000100101100100101: oled_data = 16'b1101110011010101;
				18'b000100101110100101: oled_data = 16'b1101010100110101;
				18'b000100110000100101: oled_data = 16'b1101111001011001;
				18'b000100110010100101: oled_data = 16'b1100110101010110;
				18'b000100110100100101: oled_data = 16'b1100110010010100;
				18'b000100110110100101: oled_data = 16'b1110010011010110;
				18'b000100111000100101: oled_data = 16'b1101110011010101;
				18'b000100111010100101: oled_data = 16'b1101110011010110;
				18'b000100111100100101: oled_data = 16'b1100110000110011;
				18'b000100111110100101: oled_data = 16'b1101110010010101;
				18'b000101000000100101: oled_data = 16'b1101110011010110;
				18'b000101000010100101: oled_data = 16'b1110010011010110;
				18'b000101000100100101: oled_data = 16'b1100110000010011;
				18'b000101000110100101: oled_data = 16'b1000101010101100;
				18'b000101001000100101: oled_data = 16'b0110101010001010;
				18'b000101001010100101: oled_data = 16'b0101001010001000;
				18'b000101001100100101: oled_data = 16'b0100101000100111;
				18'b000101001110100101: oled_data = 16'b0011100110000110;
				18'b000101010000100101: oled_data = 16'b0011000101000101;
				18'b000101010010100101: oled_data = 16'b0010100100000011;
				18'b000101010100100101: oled_data = 16'b0010000100000011;
				18'b000101010110100101: oled_data = 16'b0010000100000011;
				18'b000101011000100101: oled_data = 16'b0011000101100101;
				18'b000101011010100101: oled_data = 16'b0011000101000100;
				18'b000101011100100101: oled_data = 16'b0010100100100011;
				18'b000101011110100101: oled_data = 16'b0101001010001001;
				18'b000101100000100101: oled_data = 16'b1101011010111001;
				18'b000101100010100101: oled_data = 16'b1110111100111011;
				18'b000101100100100101: oled_data = 16'b1110111100011010;
				18'b000101100110100101: oled_data = 16'b1110111100011010;
				18'b000101101000100101: oled_data = 16'b1110111100011010;
				18'b000101101010100101: oled_data = 16'b1110011100011010;
				18'b000101101100100101: oled_data = 16'b1110011100011010;
				18'b000101101110100101: oled_data = 16'b1110111100011011;
				18'b000101110000100101: oled_data = 16'b1110111100011010;
				18'b000101110010100101: oled_data = 16'b1110111100011010;
				18'b000101110100100101: oled_data = 16'b1101111011011001;
				18'b000101110110100101: oled_data = 16'b1101111011011001;
				18'b000101111000100101: oled_data = 16'b1110011100011010;
				18'b000101111010100101: oled_data = 16'b1110011011011001;
				18'b000101111100100101: oled_data = 16'b1101110100110100;
				18'b000101111110100101: oled_data = 16'b1110010010110011;
				18'b000110000000100101: oled_data = 16'b1010101001101001;
				18'b000110000010100101: oled_data = 16'b1011001000101001;
				18'b000110000100100101: oled_data = 16'b1011001000101001;
				18'b000110000110100101: oled_data = 16'b1011001001001001;
				18'b000110001000100101: oled_data = 16'b1011101010101011;
				18'b000110001010100101: oled_data = 16'b1011001001101010;
				18'b000110001100100101: oled_data = 16'b1010000111100111;
				18'b000110001110100101: oled_data = 16'b1001000110100111;
				18'b000110010000100101: oled_data = 16'b1011011000011000;
				18'b000110010010100101: oled_data = 16'b1011111011111100;
				18'b000110010100100101: oled_data = 16'b1011111011111011;
				18'b000110010110100101: oled_data = 16'b1011111011111011;
				18'b000110011000100101: oled_data = 16'b1011111011111011;
				18'b000110011010100101: oled_data = 16'b1100111100111100;
				18'b000110011100100101: oled_data = 16'b1011111100011100;
				18'b000110011110100101: oled_data = 16'b1011110001010010;
				18'b000110100000100101: oled_data = 16'b1011001000001000;
				18'b000110100010100101: oled_data = 16'b1011001000101001;
				18'b000110100100100101: oled_data = 16'b1010101000101000;
				18'b000110100110100101: oled_data = 16'b1010101000101000;
				18'b000100011000100110: oled_data = 16'b0101001001100111;
				18'b000100011010100110: oled_data = 16'b1101011000001011;
				18'b000100011100100110: oled_data = 16'b1101011000101100;
				18'b000100011110100110: oled_data = 16'b1100010110101010;
				18'b000100100000100110: oled_data = 16'b1100010110001001;
				18'b000100100010100110: oled_data = 16'b1100010110001001;
				18'b000100100100100110: oled_data = 16'b1101010111101011;
				18'b000100100110100110: oled_data = 16'b1101010111101100;
				18'b000100101000100110: oled_data = 16'b1100110011101111;
				18'b000100101010100110: oled_data = 16'b1101110011010110;
				18'b000100101100100110: oled_data = 16'b1101110010110101;
				18'b000100101110100110: oled_data = 16'b1101111000111000;
				18'b000100110000100110: oled_data = 16'b1101111001010111;
				18'b000100110010100110: oled_data = 16'b1101111000011000;
				18'b000100110100100110: oled_data = 16'b1101010011110101;
				18'b000100110110100110: oled_data = 16'b1110010011010101;
				18'b000100111000100110: oled_data = 16'b1101110011010101;
				18'b000100111010100110: oled_data = 16'b1110010011010110;
				18'b000100111100100110: oled_data = 16'b1101010001110100;
				18'b000100111110100110: oled_data = 16'b1101010001010100;
				18'b000101000000100110: oled_data = 16'b1101110011010110;
				18'b000101000010100110: oled_data = 16'b1101110011010101;
				18'b000101000100100110: oled_data = 16'b1101110011010101;
				18'b000101000110100110: oled_data = 16'b1000001011101100;
				18'b000101001000100110: oled_data = 16'b0100001000000111;
				18'b000101001010100110: oled_data = 16'b0100101000100111;
				18'b000101001100100110: oled_data = 16'b0101101010101001;
				18'b000101001110100110: oled_data = 16'b0110001011101010;
				18'b000101010000100110: oled_data = 16'b0111001100101100;
				18'b000101010010100110: oled_data = 16'b1000001111101111;
				18'b000101010100100110: oled_data = 16'b1001110010110001;
				18'b000101010110100110: oled_data = 16'b1011110110110110;
				18'b000101011000100110: oled_data = 16'b0111001101001100;
				18'b000101011010100110: oled_data = 16'b0010100100100100;
				18'b000101011100100110: oled_data = 16'b0100000111100111;
				18'b000101011110100110: oled_data = 16'b1100111000111000;
				18'b000101100000100110: oled_data = 16'b1110111100111011;
				18'b000101100010100110: oled_data = 16'b1110111100011010;
				18'b000101100100100110: oled_data = 16'b1110111100011010;
				18'b000101100110100110: oled_data = 16'b1110111100011010;
				18'b000101101000100110: oled_data = 16'b1110011100011010;
				18'b000101101010100110: oled_data = 16'b1110111100011010;
				18'b000101101100100110: oled_data = 16'b1110111100011010;
				18'b000101101110100110: oled_data = 16'b1110111100011010;
				18'b000101110000100110: oled_data = 16'b1110111100011010;
				18'b000101110010100110: oled_data = 16'b1110011011111010;
				18'b000101110100100110: oled_data = 16'b1101111010111001;
				18'b000101110110100110: oled_data = 16'b1110111100011010;
				18'b000101111000100110: oled_data = 16'b1110111100111010;
				18'b000101111010100110: oled_data = 16'b1101111010011000;
				18'b000101111100100110: oled_data = 16'b1101010100010100;
				18'b000101111110100110: oled_data = 16'b1101110001110001;
				18'b000110000000100110: oled_data = 16'b1010101000101001;
				18'b000110000010100110: oled_data = 16'b1011001000101001;
				18'b000110000100100110: oled_data = 16'b1011001010001010;
				18'b000110000110100110: oled_data = 16'b1101010000110000;
				18'b000110001000100110: oled_data = 16'b1110010011110011;
				18'b000110001010100110: oled_data = 16'b1100101111001111;
				18'b000110001100100110: oled_data = 16'b1010000111101000;
				18'b000110001110100110: oled_data = 16'b1001101000101001;
				18'b000110010000100110: oled_data = 16'b1011111010111010;
				18'b000110010010100110: oled_data = 16'b1011111011111100;
				18'b000110010100100110: oled_data = 16'b1011111011111100;
				18'b000110010110100110: oled_data = 16'b1011111011111011;
				18'b000110011000100110: oled_data = 16'b1011111011111011;
				18'b000110011010100110: oled_data = 16'b1100011011111100;
				18'b000110011100100110: oled_data = 16'b1011111100011100;
				18'b000110011110100110: oled_data = 16'b1011110011110100;
				18'b000110100000100110: oled_data = 16'b1011001000001001;
				18'b000110100010100110: oled_data = 16'b1011001000101000;
				18'b000110100100100110: oled_data = 16'b1011001000101000;
				18'b000110100110100110: oled_data = 16'b1010101000101000;
				18'b000100011000100111: oled_data = 16'b0010100100000100;
				18'b000100011010100111: oled_data = 16'b0101101010000110;
				18'b000100011100100111: oled_data = 16'b1000110000101000;
				18'b000100011110100111: oled_data = 16'b1010010011101011;
				18'b000100100000100111: oled_data = 16'b1011010100101100;
				18'b000100100010100111: oled_data = 16'b1011110011101101;
				18'b000100100100100111: oled_data = 16'b1011110001001111;
				18'b000100100110100111: oled_data = 16'b1011001110001111;
				18'b000100101000100111: oled_data = 16'b1100110001010100;
				18'b000100101010100111: oled_data = 16'b1110010011010110;
				18'b000100101100100111: oled_data = 16'b1101010010110101;
				18'b000100101110100111: oled_data = 16'b1110011010011001;
				18'b000100110000100111: oled_data = 16'b1110111011111010;
				18'b000100110010100111: oled_data = 16'b1101010111010110;
				18'b000100110100100111: oled_data = 16'b1101010010110100;
				18'b000100110110100111: oled_data = 16'b1101110011010110;
				18'b000100111000100111: oled_data = 16'b1101110011010101;
				18'b000100111010100111: oled_data = 16'b1101110011010101;
				18'b000100111100100111: oled_data = 16'b1101110011010101;
				18'b000100111110100111: oled_data = 16'b1101110011010101;
				18'b000101000000100111: oled_data = 16'b1101110011010101;
				18'b000101000010100111: oled_data = 16'b1101110011010101;
				18'b000101000100100111: oled_data = 16'b1101110011010101;
				18'b000101000110100111: oled_data = 16'b1100110101010110;
				18'b000101001000100111: oled_data = 16'b1110011011011010;
				18'b000101001010100111: oled_data = 16'b1110011011111010;
				18'b000101001100100111: oled_data = 16'b1110011100011010;
				18'b000101001110100111: oled_data = 16'b1110011100011010;
				18'b000101010000100111: oled_data = 16'b1110111100011011;
				18'b000101010010100111: oled_data = 16'b1111011100111100;
				18'b000101010100100111: oled_data = 16'b1111011101111100;
				18'b000101010110100111: oled_data = 16'b1010010011010010;
				18'b000101011000100111: oled_data = 16'b0011000101000101;
				18'b000101011010100111: oled_data = 16'b0011100110000110;
				18'b000101011100100111: oled_data = 16'b1011110101110101;
				18'b000101011110100111: oled_data = 16'b1110111100111100;
				18'b000101100000100111: oled_data = 16'b1110111100011010;
				18'b000101100010100111: oled_data = 16'b1110111100011010;
				18'b000101100100100111: oled_data = 16'b1110111100011010;
				18'b000101100110100111: oled_data = 16'b1110111100011010;
				18'b000101101000100111: oled_data = 16'b1110011100011010;
				18'b000101101010100111: oled_data = 16'b1110011100011010;
				18'b000101101100100111: oled_data = 16'b1110111100011010;
				18'b000101101110100111: oled_data = 16'b1110111100011010;
				18'b000101110000100111: oled_data = 16'b1110011100011010;
				18'b000101110010100111: oled_data = 16'b1101111010011000;
				18'b000101110100100111: oled_data = 16'b1110011100011010;
				18'b000101110110100111: oled_data = 16'b1110111100111010;
				18'b000101111000100111: oled_data = 16'b1110011011111010;
				18'b000101111010100111: oled_data = 16'b1100010101010100;
				18'b000101111100100111: oled_data = 16'b1101110011110100;
				18'b000101111110100111: oled_data = 16'b1101010000110000;
				18'b000110000000100111: oled_data = 16'b1010101000101000;
				18'b000110000010100111: oled_data = 16'b1011001001001001;
				18'b000110000100100111: oled_data = 16'b1101010000110000;
				18'b000110000110100111: oled_data = 16'b1110110011110011;
				18'b000110001000100111: oled_data = 16'b1100001100101100;
				18'b000110001010100111: oled_data = 16'b1011101001001001;
				18'b000110001100100111: oled_data = 16'b1011001000101001;
				18'b000110001110100111: oled_data = 16'b1010101011101100;
				18'b000110010000100111: oled_data = 16'b1011111010111010;
				18'b000110010010100111: oled_data = 16'b1011111011011011;
				18'b000110010100100111: oled_data = 16'b1011111011111100;
				18'b000110010110100111: oled_data = 16'b1011111011111011;
				18'b000110011000100111: oled_data = 16'b1011011011011011;
				18'b000110011010100111: oled_data = 16'b1011111011011011;
				18'b000110011100100111: oled_data = 16'b1011111100011100;
				18'b000110011110100111: oled_data = 16'b1011110100110100;
				18'b000110100000100111: oled_data = 16'b1011001000001001;
				18'b000110100010100111: oled_data = 16'b1010101000001000;
				18'b000110100100100111: oled_data = 16'b1010100111101000;
				18'b000110100110100111: oled_data = 16'b1010101000001000;
				18'b000100011000101000: oled_data = 16'b0011100110100100;
				18'b000100011010101000: oled_data = 16'b0100101000100110;
				18'b000100011100101000: oled_data = 16'b0101101011001000;
				18'b000100011110101000: oled_data = 16'b0110101101001100;
				18'b000100100000101000: oled_data = 16'b1000110000010000;
				18'b000100100010101000: oled_data = 16'b1010101110110001;
				18'b000100100100101000: oled_data = 16'b1011001101010001;
				18'b000100100110101000: oled_data = 16'b1011001101110001;
				18'b000100101000101000: oled_data = 16'b1101110010110101;
				18'b000100101010101000: oled_data = 16'b1110010011010110;
				18'b000100101100101000: oled_data = 16'b1101010010110101;
				18'b000100101110101000: oled_data = 16'b1110011010011001;
				18'b000100110000101000: oled_data = 16'b1110111100011010;
				18'b000100110010101000: oled_data = 16'b1110011010111001;
				18'b000100110100101000: oled_data = 16'b1101010011110101;
				18'b000100110110101000: oled_data = 16'b1101110011010101;
				18'b000100111000101000: oled_data = 16'b1101110011010101;
				18'b000100111010101000: oled_data = 16'b1101110011010101;
				18'b000100111100101000: oled_data = 16'b1101110011010101;
				18'b000100111110101000: oled_data = 16'b1101110011010101;
				18'b000101000000101000: oled_data = 16'b1101110011010101;
				18'b000101000010101000: oled_data = 16'b1101110011010101;
				18'b000101000100101000: oled_data = 16'b1101110010110101;
				18'b000101000110101000: oled_data = 16'b1101010100110110;
				18'b000101001000101000: oled_data = 16'b1110111100011011;
				18'b000101001010101000: oled_data = 16'b1110111100011010;
				18'b000101001100101000: oled_data = 16'b1110111100011010;
				18'b000101001110101000: oled_data = 16'b1110011100011010;
				18'b000101010000101000: oled_data = 16'b1110011100011010;
				18'b000101010010101000: oled_data = 16'b1111011100111100;
				18'b000101010100101000: oled_data = 16'b1010110011110011;
				18'b000101010110101000: oled_data = 16'b0011000101000101;
				18'b000101011000101000: oled_data = 16'b0011100110000110;
				18'b000101011010101000: oled_data = 16'b1011010101010100;
				18'b000101011100101000: oled_data = 16'b1110111101011100;
				18'b000101011110101000: oled_data = 16'b1110011100011010;
				18'b000101100000101000: oled_data = 16'b1110111100011010;
				18'b000101100010101000: oled_data = 16'b1110111100011010;
				18'b000101100100101000: oled_data = 16'b1110111100011010;
				18'b000101100110101000: oled_data = 16'b1110111100011010;
				18'b000101101000101000: oled_data = 16'b1110011100011010;
				18'b000101101010101000: oled_data = 16'b1110111100011010;
				18'b000101101100101000: oled_data = 16'b1110111100011010;
				18'b000101101110101000: oled_data = 16'b1110111100011010;
				18'b000101110000101000: oled_data = 16'b1101111010011000;
				18'b000101110010101000: oled_data = 16'b1110011011111010;
				18'b000101110100101000: oled_data = 16'b1110111100111010;
				18'b000101110110101000: oled_data = 16'b1101111011011001;
				18'b000101111000101000: oled_data = 16'b1100110101010101;
				18'b000101111010101000: oled_data = 16'b1101010110010101;
				18'b000101111100101000: oled_data = 16'b1110010100010100;
				18'b000101111110101000: oled_data = 16'b1101001111001111;
				18'b000110000000101000: oled_data = 16'b1010101000001000;
				18'b000110000010101000: oled_data = 16'b1100001011101100;
				18'b000110000100101000: oled_data = 16'b1110110011110011;
				18'b000110000110101000: oled_data = 16'b1100101101101110;
				18'b000110001000101000: oled_data = 16'b1011001000101001;
				18'b000110001010101000: oled_data = 16'b1011001001001001;
				18'b000110001100101000: oled_data = 16'b1011001000101001;
				18'b000110001110101000: oled_data = 16'b1011001011101100;
				18'b000110010000101000: oled_data = 16'b1011111010111010;
				18'b000110010010101000: oled_data = 16'b1011111011111100;
				18'b000110010100101000: oled_data = 16'b1011111011011011;
				18'b000110010110101000: oled_data = 16'b1010011000111001;
				18'b000110011000101000: oled_data = 16'b1001010111011000;
				18'b000110011010101000: oled_data = 16'b1010111001111010;
				18'b000110011100101000: oled_data = 16'b1011111100011100;
				18'b000110011110101000: oled_data = 16'b1011010100010100;
				18'b000110100000101000: oled_data = 16'b1010100111101000;
				18'b000110100010101000: oled_data = 16'b1010001000001000;
				18'b000110100100101000: oled_data = 16'b1010101000001000;
				18'b000110100110101000: oled_data = 16'b1010101000001000;
				18'b000100011000101001: oled_data = 16'b0111101111101001;
				18'b000100011010101001: oled_data = 16'b0111101111001010;
				18'b000100011100101001: oled_data = 16'b1000001111101011;
				18'b000100011110101001: oled_data = 16'b0110101101001011;
				18'b000100100000101001: oled_data = 16'b0110101010101011;
				18'b000100100010101001: oled_data = 16'b1011001110110001;
				18'b000100100100101001: oled_data = 16'b1010101100110000;
				18'b000100100110101001: oled_data = 16'b1101010001010100;
				18'b000100101000101001: oled_data = 16'b1110010011010110;
				18'b000100101010101001: oled_data = 16'b1101110011010101;
				18'b000100101100101001: oled_data = 16'b1101110011010101;
				18'b000100101110101001: oled_data = 16'b1101111001111000;
				18'b000100110000101001: oled_data = 16'b1110111100011010;
				18'b000100110010101001: oled_data = 16'b1110011011011001;
				18'b000100110100101001: oled_data = 16'b1101010100010101;
				18'b000100110110101001: oled_data = 16'b1101110011010101;
				18'b000100111000101001: oled_data = 16'b1101110011010101;
				18'b000100111010101001: oled_data = 16'b1101110011010101;
				18'b000100111100101001: oled_data = 16'b1101110011010101;
				18'b000100111110101001: oled_data = 16'b1101110011010101;
				18'b000101000000101001: oled_data = 16'b1101110011010101;
				18'b000101000010101001: oled_data = 16'b1101110011010101;
				18'b000101000100101001: oled_data = 16'b1101110010110101;
				18'b000101000110101001: oled_data = 16'b1101110101010110;
				18'b000101001000101001: oled_data = 16'b1110111011111010;
				18'b000101001010101001: oled_data = 16'b1110111100011010;
				18'b000101001100101001: oled_data = 16'b1110111100011010;
				18'b000101001110101001: oled_data = 16'b1110111100011010;
				18'b000101010000101001: oled_data = 16'b1111011101011011;
				18'b000101010010101001: oled_data = 16'b1010110100110011;
				18'b000101010100101001: oled_data = 16'b0011100101100101;
				18'b000101010110101001: oled_data = 16'b0011100101100101;
				18'b000101011000101001: oled_data = 16'b1010110100110100;
				18'b000101011010101001: oled_data = 16'b1110111100111011;
				18'b000101011100101001: oled_data = 16'b1110011100011010;
				18'b000101011110101001: oled_data = 16'b1110011100011010;
				18'b000101100000101001: oled_data = 16'b1110011100011010;
				18'b000101100010101001: oled_data = 16'b1110011100011010;
				18'b000101100100101001: oled_data = 16'b1110111100011010;
				18'b000101100110101001: oled_data = 16'b1110111100011010;
				18'b000101101000101001: oled_data = 16'b1110111100011010;
				18'b000101101010101001: oled_data = 16'b1110111100011010;
				18'b000101101100101001: oled_data = 16'b1110111100011010;
				18'b000101101110101001: oled_data = 16'b1101111010111001;
				18'b000101110000101001: oled_data = 16'b1101111011011001;
				18'b000101110010101001: oled_data = 16'b1110111100111011;
				18'b000101110100101001: oled_data = 16'b1110011011111010;
				18'b000101110110101001: oled_data = 16'b1100010100110100;
				18'b000101111000101001: oled_data = 16'b1100110101110101;
				18'b000101111010101001: oled_data = 16'b1110111010011001;
				18'b000101111100101001: oled_data = 16'b1110010100110100;
				18'b000101111110101001: oled_data = 16'b1100101110001110;
				18'b000110000000101001: oled_data = 16'b1011001000001000;
				18'b000110000010101001: oled_data = 16'b1100101110101110;
				18'b000110000100101001: oled_data = 16'b1110010011010010;
				18'b000110000110101001: oled_data = 16'b1011101010001010;
				18'b000110001000101001: oled_data = 16'b1011101000101001;
				18'b000110001010101001: oled_data = 16'b1011101001001001;
				18'b000110001100101001: oled_data = 16'b1011001000101001;
				18'b000110001110101001: oled_data = 16'b1011001010101011;
				18'b000110010000101001: oled_data = 16'b1011111001111001;
				18'b000110010010101001: oled_data = 16'b1011111011111100;
				18'b000110010100101001: oled_data = 16'b1010111001011001;
				18'b000110010110101001: oled_data = 16'b1001010110111000;
				18'b000110011000101001: oled_data = 16'b1001010111011000;
				18'b000110011010101001: oled_data = 16'b1010011000011001;
				18'b000110011100101001: oled_data = 16'b1010111010111011;
				18'b000110011110101001: oled_data = 16'b1010010001010001;
				18'b000110100000101001: oled_data = 16'b1010100111101000;
				18'b000110100010101001: oled_data = 16'b1010101000101001;
				18'b000110100100101001: oled_data = 16'b1010101000101001;
				18'b000110100110101001: oled_data = 16'b1011001000001000;
				18'b000100011000101010: oled_data = 16'b0111101111001011;
				18'b000100011010101010: oled_data = 16'b0101101010100111;
				18'b000100011100101010: oled_data = 16'b0111001101101001;
				18'b000100011110101010: oled_data = 16'b0110101101001100;
				18'b000100100000101010: oled_data = 16'b1010001110110001;
				18'b000100100010101010: oled_data = 16'b1011101110010001;
				18'b000100100100101010: oled_data = 16'b1100001111010010;
				18'b000100100110101010: oled_data = 16'b1101110011010101;
				18'b000100101000101010: oled_data = 16'b1101110011010101;
				18'b000100101010101010: oled_data = 16'b1101110011010101;
				18'b000100101100101010: oled_data = 16'b1101110011010101;
				18'b000100101110101010: oled_data = 16'b1101110110110111;
				18'b000100110000101010: oled_data = 16'b1110111100011011;
				18'b000100110010101010: oled_data = 16'b1110011011011010;
				18'b000100110100101010: oled_data = 16'b1101010100010101;
				18'b000100110110101010: oled_data = 16'b1101110011010110;
				18'b000100111000101010: oled_data = 16'b1101110011010101;
				18'b000100111010101010: oled_data = 16'b1101110011010101;
				18'b000100111100101010: oled_data = 16'b1101110011010101;
				18'b000100111110101010: oled_data = 16'b1101110011010101;
				18'b000101000000101010: oled_data = 16'b1101110011010101;
				18'b000101000010101010: oled_data = 16'b1101110011010101;
				18'b000101000100101010: oled_data = 16'b1101110010110101;
				18'b000101000110101010: oled_data = 16'b1101110101010110;
				18'b000101001000101010: oled_data = 16'b1110011011111010;
				18'b000101001010101010: oled_data = 16'b1110111100011010;
				18'b000101001100101010: oled_data = 16'b1110111100011010;
				18'b000101001110101010: oled_data = 16'b1110111101011011;
				18'b000101010000101010: oled_data = 16'b1010110100110011;
				18'b000101010010101010: oled_data = 16'b0011100110000110;
				18'b000101010100101010: oled_data = 16'b0100000111000110;
				18'b000101010110101010: oled_data = 16'b1011010101010101;
				18'b000101011000101010: oled_data = 16'b1111011101011100;
				18'b000101011010101010: oled_data = 16'b1110111100011010;
				18'b000101011100101010: oled_data = 16'b1110111100011010;
				18'b000101011110101010: oled_data = 16'b1110111100011010;
				18'b000101100000101010: oled_data = 16'b1110111100011010;
				18'b000101100010101010: oled_data = 16'b1110111100011010;
				18'b000101100100101010: oled_data = 16'b1110111100011010;
				18'b000101100110101010: oled_data = 16'b1110111100011010;
				18'b000101101000101010: oled_data = 16'b1110111100011010;
				18'b000101101010101010: oled_data = 16'b1110111100011010;
				18'b000101101100101010: oled_data = 16'b1110111100011010;
				18'b000101101110101010: oled_data = 16'b1110011011111010;
				18'b000101110000101010: oled_data = 16'b1110111100111011;
				18'b000101110010101010: oled_data = 16'b1110011010011001;
				18'b000101110100101010: oled_data = 16'b1101010101010101;
				18'b000101110110101010: oled_data = 16'b1101110101110110;
				18'b000101111000101010: oled_data = 16'b1110111011011010;
				18'b000101111010101010: oled_data = 16'b1110011011011010;
				18'b000101111100101010: oled_data = 16'b1101110100110100;
				18'b000101111110101010: oled_data = 16'b1100001101001101;
				18'b000110000000101010: oled_data = 16'b1011001000101001;
				18'b000110000010101010: oled_data = 16'b1101010000110000;
				18'b000110000100101010: oled_data = 16'b1101010000010000;
				18'b000110000110101010: oled_data = 16'b1011001001001001;
				18'b000110001000101010: oled_data = 16'b1011101001001001;
				18'b000110001010101010: oled_data = 16'b1011001001001001;
				18'b000110001100101010: oled_data = 16'b1011001001001001;
				18'b000110001110101010: oled_data = 16'b1011001000101001;
				18'b000110010000101010: oled_data = 16'b1011110101010101;
				18'b000110010010101010: oled_data = 16'b1011111100011100;
				18'b000110010100101010: oled_data = 16'b1001111000011000;
				18'b000110010110101010: oled_data = 16'b1001010111011000;
				18'b000110011000101010: oled_data = 16'b1001010111011000;
				18'b000110011010101010: oled_data = 16'b1001010111011000;
				18'b000110011100101010: oled_data = 16'b1010111001011000;
				18'b000110011110101010: oled_data = 16'b1010101011101100;
				18'b000110100000101010: oled_data = 16'b1010101000001000;
				18'b000110100010101010: oled_data = 16'b1010101000101000;
				18'b000110100100101010: oled_data = 16'b1010101000001000;
				18'b000110100110101010: oled_data = 16'b1010101000001000;
				18'b000100011000101011: oled_data = 16'b0111101110101011;
				18'b000100011010101011: oled_data = 16'b0111001110001011;
				18'b000100011100101011: oled_data = 16'b1000010000001100;
				18'b000100011110101011: oled_data = 16'b1001010000001111;
				18'b000100100000101011: oled_data = 16'b1101010010010101;
				18'b000100100010101011: oled_data = 16'b1100110001010100;
				18'b000100100100101011: oled_data = 16'b1101110011010110;
				18'b000100100110101011: oled_data = 16'b1101110011010101;
				18'b000100101000101011: oled_data = 16'b1101110011010101;
				18'b000100101010101011: oled_data = 16'b1101110011010101;
				18'b000100101100101011: oled_data = 16'b1101110011010101;
				18'b000100101110101011: oled_data = 16'b1100010010010011;
				18'b000100110000101011: oled_data = 16'b1110111011111010;
				18'b000100110010101011: oled_data = 16'b1110011011111010;
				18'b000100110100101011: oled_data = 16'b1101010100010101;
				18'b000100110110101011: oled_data = 16'b1101110011010110;
				18'b000100111000101011: oled_data = 16'b1101110011010101;
				18'b000100111010101011: oled_data = 16'b1101110011010101;
				18'b000100111100101011: oled_data = 16'b1101110011010101;
				18'b000100111110101011: oled_data = 16'b1101110011010101;
				18'b000101000000101011: oled_data = 16'b1101110011010101;
				18'b000101000010101011: oled_data = 16'b1101110011010101;
				18'b000101000100101011: oled_data = 16'b1101110010110101;
				18'b000101000110101011: oled_data = 16'b1101110101010110;
				18'b000101001000101011: oled_data = 16'b1110011011111010;
				18'b000101001010101011: oled_data = 16'b1110111100011010;
				18'b000101001100101011: oled_data = 16'b1110111101011011;
				18'b000101001110101011: oled_data = 16'b1011010110010100;
				18'b000101010000101011: oled_data = 16'b0011000101000100;
				18'b000101010010101011: oled_data = 16'b0101001000101000;
				18'b000101010100101011: oled_data = 16'b1100110111110111;
				18'b000101010110101011: oled_data = 16'b1110111100111100;
				18'b000101011000101011: oled_data = 16'b1110111100011011;
				18'b000101011010101011: oled_data = 16'b1110111100011011;
				18'b000101011100101011: oled_data = 16'b1110111100011010;
				18'b000101011110101011: oled_data = 16'b1110111100011010;
				18'b000101100000101011: oled_data = 16'b1110111100011010;
				18'b000101100010101011: oled_data = 16'b1110111100011010;
				18'b000101100100101011: oled_data = 16'b1110111100011010;
				18'b000101100110101011: oled_data = 16'b1110111100011010;
				18'b000101101000101011: oled_data = 16'b1110111100011010;
				18'b000101101010101011: oled_data = 16'b1110111100011010;
				18'b000101101100101011: oled_data = 16'b1110111100011011;
				18'b000101101110101011: oled_data = 16'b1110111100111011;
				18'b000101110000101011: oled_data = 16'b1101011001111000;
				18'b000101110010101011: oled_data = 16'b1100110100110100;
				18'b000101110100101011: oled_data = 16'b1101110101010101;
				18'b000101110110101011: oled_data = 16'b1110111010111001;
				18'b000101111000101011: oled_data = 16'b1110111100011011;
				18'b000101111010101011: oled_data = 16'b1110011011011010;
				18'b000101111100101011: oled_data = 16'b1101110101010100;
				18'b000101111110101011: oled_data = 16'b1011101100001100;
				18'b000110000000101011: oled_data = 16'b1011001000101001;
				18'b000110000010101011: oled_data = 16'b1101110001110001;
				18'b000110000100101011: oled_data = 16'b1100101101101101;
				18'b000110000110101011: oled_data = 16'b1011001000101001;
				18'b000110001000101011: oled_data = 16'b1011001001001001;
				18'b000110001010101011: oled_data = 16'b1011001001001001;
				18'b000110001100101011: oled_data = 16'b1011001001001001;
				18'b000110001110101011: oled_data = 16'b1011001000101001;
				18'b000110010000101011: oled_data = 16'b1010101011101011;
				18'b000110010010101011: oled_data = 16'b1011111010111010;
				18'b000110010100101011: oled_data = 16'b1010011001011010;
				18'b000110010110101011: oled_data = 16'b1000110111011000;
				18'b000110011000101011: oled_data = 16'b1001010111111001;
				18'b000110011010101011: oled_data = 16'b1001111000011001;
				18'b000110011100101011: oled_data = 16'b1011010001110010;
				18'b000110011110101011: oled_data = 16'b1011001000101001;
				18'b000110100000101011: oled_data = 16'b1010101000101001;
				18'b000110100010101011: oled_data = 16'b1010101000001000;
				18'b000110100100101011: oled_data = 16'b1010101000001000;
				18'b000110100110101011: oled_data = 16'b1010101000001000;
				18'b000100011000101100: oled_data = 16'b1000110001101110;
				18'b000100011010101100: oled_data = 16'b1000110001101111;
				18'b000100011100101100: oled_data = 16'b1000001111001101;
				18'b000100011110101100: oled_data = 16'b1011110010010011;
				18'b000100100000101100: oled_data = 16'b1101010001110100;
				18'b000100100010101100: oled_data = 16'b1101110010110101;
				18'b000100100100101100: oled_data = 16'b1101110011010101;
				18'b000100100110101100: oled_data = 16'b1101110011010101;
				18'b000100101000101100: oled_data = 16'b1101110011010101;
				18'b000100101010101100: oled_data = 16'b1101110011010110;
				18'b000100101100101100: oled_data = 16'b1101110010010101;
				18'b000100101110101100: oled_data = 16'b1011001110010001;
				18'b000100110000101100: oled_data = 16'b1100110101110110;
				18'b000100110010101100: oled_data = 16'b1110111011111010;
				18'b000100110100101100: oled_data = 16'b1101010011110101;
				18'b000100110110101100: oled_data = 16'b1101110011010101;
				18'b000100111000101100: oled_data = 16'b1101110011010101;
				18'b000100111010101100: oled_data = 16'b1101110011010101;
				18'b000100111100101100: oled_data = 16'b1101110011010101;
				18'b000100111110101100: oled_data = 16'b1101110011010101;
				18'b000101000000101100: oled_data = 16'b1101110011010101;
				18'b000101000010101100: oled_data = 16'b1101110011010101;
				18'b000101000100101100: oled_data = 16'b1101110010110101;
				18'b000101000110101100: oled_data = 16'b1101010101010110;
				18'b000101001000101100: oled_data = 16'b1110111011111010;
				18'b000101001010101100: oled_data = 16'b1110111100011010;
				18'b000101001100101100: oled_data = 16'b1101111011011001;
				18'b000101001110101100: oled_data = 16'b0101001001000111;
				18'b000101010000101100: oled_data = 16'b0110001011001001;
				18'b000101010010101100: oled_data = 16'b1101011001111000;
				18'b000101010100101100: oled_data = 16'b1110111100111011;
				18'b000101010110101100: oled_data = 16'b1110111100011011;
				18'b000101011000101100: oled_data = 16'b1110111100011011;
				18'b000101011010101100: oled_data = 16'b1110111100011010;
				18'b000101011100101100: oled_data = 16'b1110111100011010;
				18'b000101011110101100: oled_data = 16'b1110111100011010;
				18'b000101100000101100: oled_data = 16'b1110111100011010;
				18'b000101100010101100: oled_data = 16'b1110111100011010;
				18'b000101100100101100: oled_data = 16'b1110111100011010;
				18'b000101100110101100: oled_data = 16'b1110111100011010;
				18'b000101101000101100: oled_data = 16'b1110111100011010;
				18'b000101101010101100: oled_data = 16'b1110111100111011;
				18'b000101101100101100: oled_data = 16'b1110011011111010;
				18'b000101101110101100: oled_data = 16'b1101010110010110;
				18'b000101110000101100: oled_data = 16'b1100110100110100;
				18'b000101110010101100: oled_data = 16'b1101110100110101;
				18'b000101110100101100: oled_data = 16'b1110011000011000;
				18'b000101110110101100: oled_data = 16'b1110111100011010;
				18'b000101111000101100: oled_data = 16'b1110011100011010;
				18'b000101111010101100: oled_data = 16'b1110111100011010;
				18'b000101111100101100: oled_data = 16'b1101010101110101;
				18'b000101111110101100: oled_data = 16'b1011101011101100;
				18'b000110000000101100: oled_data = 16'b1011001001001001;
				18'b000110000010101100: oled_data = 16'b1101110010010010;
				18'b000110000100101100: oled_data = 16'b1100001011101100;
				18'b000110000110101100: oled_data = 16'b1011001000101001;
				18'b000110001000101100: oled_data = 16'b1011001001001001;
				18'b000110001010101100: oled_data = 16'b1011001001001001;
				18'b000110001100101100: oled_data = 16'b1011001001001001;
				18'b000110001110101100: oled_data = 16'b1011101001001001;
				18'b000110010000101100: oled_data = 16'b1001100110100111;
				18'b000110010010101100: oled_data = 16'b1001101010101011;
				18'b000110010100101100: oled_data = 16'b1011110100110101;
				18'b000110010110101100: oled_data = 16'b1010010101110110;
				18'b000110011000101100: oled_data = 16'b1010010100110101;
				18'b000110011010101100: oled_data = 16'b1010110000010001;
				18'b000110011100101100: oled_data = 16'b1011001001001001;
				18'b000110011110101100: oled_data = 16'b1011001000101001;
				18'b000110100000101100: oled_data = 16'b1011001000101000;
				18'b000110100010101100: oled_data = 16'b1010101000001000;
				18'b000110100100101100: oled_data = 16'b1010101000001000;
				18'b000110100110101100: oled_data = 16'b1010101000001000;
				18'b000100011000101101: oled_data = 16'b0101101011101010;
				18'b000100011010101101: oled_data = 16'b0100001000100111;
				18'b000100011100101101: oled_data = 16'b1000101101001110;
				18'b000100011110101101: oled_data = 16'b1101010010010101;
				18'b000100100000101101: oled_data = 16'b1101110010110101;
				18'b000100100010101101: oled_data = 16'b1101110011010101;
				18'b000100100100101101: oled_data = 16'b1101110011010101;
				18'b000100100110101101: oled_data = 16'b1101110011010101;
				18'b000100101000101101: oled_data = 16'b1101110011010101;
				18'b000100101010101101: oled_data = 16'b1101110011010110;
				18'b000100101100101101: oled_data = 16'b1101010001010100;
				18'b000100101110101101: oled_data = 16'b1011101101110001;
				18'b000100110000101101: oled_data = 16'b1011001110110001;
				18'b000100110010101101: oled_data = 16'b1101010111010111;
				18'b000100110100101101: oled_data = 16'b1101110100010110;
				18'b000100110110101101: oled_data = 16'b1101110011010101;
				18'b000100111000101101: oled_data = 16'b1101110011010101;
				18'b000100111010101101: oled_data = 16'b1101110011010101;
				18'b000100111100101101: oled_data = 16'b1101110011010101;
				18'b000100111110101101: oled_data = 16'b1101110011010101;
				18'b000101000000101101: oled_data = 16'b1101110011010101;
				18'b000101000010101101: oled_data = 16'b1101110010110101;
				18'b000101000100101101: oled_data = 16'b1101110010110101;
				18'b000101000110101101: oled_data = 16'b1101010101010110;
				18'b000101001000101101: oled_data = 16'b1110111100011010;
				18'b000101001010101101: oled_data = 16'b1110111100111011;
				18'b000101001100101101: oled_data = 16'b1011010101010100;
				18'b000101001110101101: oled_data = 16'b0111001101101100;
				18'b000101010000101101: oled_data = 16'b1101111011011001;
				18'b000101010010101101: oled_data = 16'b1110111100111011;
				18'b000101010100101101: oled_data = 16'b1110111100011010;
				18'b000101010110101101: oled_data = 16'b1110111100011010;
				18'b000101011000101101: oled_data = 16'b1110111100011010;
				18'b000101011010101101: oled_data = 16'b1110111100011010;
				18'b000101011100101101: oled_data = 16'b1110111100011010;
				18'b000101011110101101: oled_data = 16'b1110111100011010;
				18'b000101100000101101: oled_data = 16'b1110111100011010;
				18'b000101100010101101: oled_data = 16'b1110111100011010;
				18'b000101100100101101: oled_data = 16'b1110111100011010;
				18'b000101100110101101: oled_data = 16'b1110111100111011;
				18'b000101101000101101: oled_data = 16'b1110111100011011;
				18'b000101101010101101: oled_data = 16'b1101111000110111;
				18'b000101101100101101: oled_data = 16'b1011010001010001;
				18'b000101101110101101: oled_data = 16'b1100110010010011;
				18'b000101110000101101: oled_data = 16'b1101110101010101;
				18'b000101110010101101: oled_data = 16'b1101010101010101;
				18'b000101110100101101: oled_data = 16'b1110011010011001;
				18'b000101110110101101: oled_data = 16'b1110011100011010;
				18'b000101111000101101: oled_data = 16'b1110011100011010;
				18'b000101111010101101: oled_data = 16'b1110111100011010;
				18'b000101111100101101: oled_data = 16'b1101010110110110;
				18'b000101111110101101: oled_data = 16'b1011101011001100;
				18'b000110000000101101: oled_data = 16'b1011001001001001;
				18'b000110000010101101: oled_data = 16'b1101010001110001;
				18'b000110000100101101: oled_data = 16'b1011101010101011;
				18'b000110000110101101: oled_data = 16'b1011001000101001;
				18'b000110001000101101: oled_data = 16'b1011001001001001;
				18'b000110001010101101: oled_data = 16'b1011001001001001;
				18'b000110001100101101: oled_data = 16'b1011001001001001;
				18'b000110001110101101: oled_data = 16'b1011101001001001;
				18'b000110010000101101: oled_data = 16'b1001100111101000;
				18'b000110010010101101: oled_data = 16'b1000000101000101;
				18'b000110010100101101: oled_data = 16'b1001100110100111;
				18'b000110010110101101: oled_data = 16'b1010101001101001;
				18'b000110011000101101: oled_data = 16'b1010101001001001;
				18'b000110011010101101: oled_data = 16'b1011001000001001;
				18'b000110011100101101: oled_data = 16'b1011001000101001;
				18'b000110011110101101: oled_data = 16'b1011001000101000;
				18'b000110100000101101: oled_data = 16'b1011001000001000;
				18'b000110100010101101: oled_data = 16'b1010101000001000;
				18'b000110100100101101: oled_data = 16'b1010101000001000;
				18'b000110100110101101: oled_data = 16'b1010101000001000;
				18'b000100011000101110: oled_data = 16'b0010100110100110;
				18'b000100011010101110: oled_data = 16'b0110001010001010;
				18'b000100011100101110: oled_data = 16'b1101010001110100;
				18'b000100011110101110: oled_data = 16'b1101110010010101;
				18'b000100100000101110: oled_data = 16'b1101110010110101;
				18'b000100100010101110: oled_data = 16'b1101110010110101;
				18'b000100100100101110: oled_data = 16'b1101110010110101;
				18'b000100100110101110: oled_data = 16'b1101110010110101;
				18'b000100101000101110: oled_data = 16'b1101110010110101;
				18'b000100101010101110: oled_data = 16'b1101110010110101;
				18'b000100101100101110: oled_data = 16'b1100001111110010;
				18'b000100101110101110: oled_data = 16'b1011001101110000;
				18'b000100110000101110: oled_data = 16'b1011001101110001;
				18'b000100110010101110: oled_data = 16'b1011001110010001;
				18'b000100110100101110: oled_data = 16'b1101010001110100;
				18'b000100110110101110: oled_data = 16'b1101110011010101;
				18'b000100111000101110: oled_data = 16'b1101110010110101;
				18'b000100111010101110: oled_data = 16'b1101110010110101;
				18'b000100111100101110: oled_data = 16'b1101110010110101;
				18'b000100111110101110: oled_data = 16'b1101110010110101;
				18'b000101000000101110: oled_data = 16'b1101110011010101;
				18'b000101000010101110: oled_data = 16'b1101110010110101;
				18'b000101000100101110: oled_data = 16'b1101110010110101;
				18'b000101000110101110: oled_data = 16'b1101010101010110;
				18'b000101001000101110: oled_data = 16'b1110111100011011;
				18'b000101001010101110: oled_data = 16'b1110111100011010;
				18'b000101001100101110: oled_data = 16'b1110011011111010;
				18'b000101001110101110: oled_data = 16'b1110011100011010;
				18'b000101010000101110: oled_data = 16'b1110011100011010;
				18'b000101010010101110: oled_data = 16'b1110011100011010;
				18'b000101010100101110: oled_data = 16'b1110111100011010;
				18'b000101010110101110: oled_data = 16'b1110011100011010;
				18'b000101011000101110: oled_data = 16'b1110011100011010;
				18'b000101011010101110: oled_data = 16'b1110011100011010;
				18'b000101011100101110: oled_data = 16'b1110111100011010;
				18'b000101011110101110: oled_data = 16'b1110111100011010;
				18'b000101100000101110: oled_data = 16'b1110111100011010;
				18'b000101100010101110: oled_data = 16'b1110111100111011;
				18'b000101100100101110: oled_data = 16'b1110111100111011;
				18'b000101100110101110: oled_data = 16'b1101111001011000;
				18'b000101101000101110: oled_data = 16'b1100010011110011;
				18'b000101101010101110: oled_data = 16'b1011001111010000;
				18'b000101101100101110: oled_data = 16'b1011110000010001;
				18'b000101101110101110: oled_data = 16'b1110010101010110;
				18'b000101110000101110: oled_data = 16'b1110010100110101;
				18'b000101110010101110: oled_data = 16'b1101010100110101;
				18'b000101110100101110: oled_data = 16'b1110011010111010;
				18'b000101110110101110: oled_data = 16'b1110011100011010;
				18'b000101111000101110: oled_data = 16'b1110011011111010;
				18'b000101111010101110: oled_data = 16'b1110111100011010;
				18'b000101111100101110: oled_data = 16'b1101111000110111;
				18'b000101111110101110: oled_data = 16'b1011001011001100;
				18'b000110000000101110: oled_data = 16'b1011001001101010;
				18'b000110000010101110: oled_data = 16'b1101010000110000;
				18'b000110000100101110: oled_data = 16'b1011101001101010;
				18'b000110000110101110: oled_data = 16'b1011101000101001;
				18'b000110001000101110: oled_data = 16'b1011001001001001;
				18'b000110001010101110: oled_data = 16'b1011001000101001;
				18'b000110001100101110: oled_data = 16'b1011001000101001;
				18'b000110001110101110: oled_data = 16'b1011001001001001;
				18'b000110010000101110: oled_data = 16'b1001100111001000;
				18'b000110010010101110: oled_data = 16'b1000000101000110;
				18'b000110010100101110: oled_data = 16'b1000000100100101;
				18'b000110010110101110: oled_data = 16'b1001100111000111;
				18'b000110011000101110: oled_data = 16'b1010101000101000;
				18'b000110011010101110: oled_data = 16'b1010000111101000;
				18'b000110011100101110: oled_data = 16'b1010101000001000;
				18'b000110011110101110: oled_data = 16'b1010101000001000;
				18'b000110100000101110: oled_data = 16'b1011001000001000;
				18'b000110100010101110: oled_data = 16'b1010101000001000;
				18'b000110100100101110: oled_data = 16'b1010100111101000;
				18'b000110100110101110: oled_data = 16'b1010100111101000;
				18'b000100011000101111: oled_data = 16'b0101001000101000;
				18'b000100011010101111: oled_data = 16'b1011010000010010;
				18'b000100011100101111: oled_data = 16'b1101010001110100;
				18'b000100011110101111: oled_data = 16'b1101110010110101;
				18'b000100100000101111: oled_data = 16'b1101110010110101;
				18'b000100100010101111: oled_data = 16'b1101110010110101;
				18'b000100100100101111: oled_data = 16'b1101110010010101;
				18'b000100100110101111: oled_data = 16'b1101110010010101;
				18'b000100101000101111: oled_data = 16'b1101110010110101;
				18'b000100101010101111: oled_data = 16'b1101010010010100;
				18'b000100101100101111: oled_data = 16'b1011001110010001;
				18'b000100101110101111: oled_data = 16'b1011001101010000;
				18'b000100110000101111: oled_data = 16'b1011001101110001;
				18'b000100110010101111: oled_data = 16'b1011001101010000;
				18'b000100110100101111: oled_data = 16'b1101010001010100;
				18'b000100110110101111: oled_data = 16'b1101110010110101;
				18'b000100111000101111: oled_data = 16'b1101110010110101;
				18'b000100111010101111: oled_data = 16'b1101110010110101;
				18'b000100111100101111: oled_data = 16'b1101110010110101;
				18'b000100111110101111: oled_data = 16'b1101110010110101;
				18'b000101000000101111: oled_data = 16'b1101110010110101;
				18'b000101000010101111: oled_data = 16'b1101110010110101;
				18'b000101000100101111: oled_data = 16'b1101110010010101;
				18'b000101000110101111: oled_data = 16'b1101010110010111;
				18'b000101001000101111: oled_data = 16'b1110011100011011;
				18'b000101001010101111: oled_data = 16'b1110011011111010;
				18'b000101001100101111: oled_data = 16'b1110011100011010;
				18'b000101001110101111: oled_data = 16'b1110011100011010;
				18'b000101010000101111: oled_data = 16'b1110011011111010;
				18'b000101010010101111: oled_data = 16'b1110011011111010;
				18'b000101010100101111: oled_data = 16'b1110011011111010;
				18'b000101010110101111: oled_data = 16'b1110011011111010;
				18'b000101011000101111: oled_data = 16'b1110011100011010;
				18'b000101011010101111: oled_data = 16'b1110011100011010;
				18'b000101011100101111: oled_data = 16'b1110111100111010;
				18'b000101011110101111: oled_data = 16'b1110111100111010;
				18'b000101100000101111: oled_data = 16'b1101111011011001;
				18'b000101100010101111: oled_data = 16'b1100110111010110;
				18'b000101100100101111: oled_data = 16'b1011110010010010;
				18'b000101100110101111: oled_data = 16'b1011001111110000;
				18'b000101101000101111: oled_data = 16'b1011101111010000;
				18'b000101101010101111: oled_data = 16'b1011101111010000;
				18'b000101101100101111: oled_data = 16'b1101110011110100;
				18'b000101101110101111: oled_data = 16'b1110010101010110;
				18'b000101110000101111: oled_data = 16'b1101110100110101;
				18'b000101110010101111: oled_data = 16'b1101010101010101;
				18'b000101110100101111: oled_data = 16'b1110011011011010;
				18'b000101110110101111: oled_data = 16'b1110011011111010;
				18'b000101111000101111: oled_data = 16'b1110011011111010;
				18'b000101111010101111: oled_data = 16'b1110011100011010;
				18'b000101111100101111: oled_data = 16'b1110011011011001;
				18'b000101111110101111: oled_data = 16'b1011001100001100;
				18'b000110000000101111: oled_data = 16'b1011001001101010;
				18'b000110000010101111: oled_data = 16'b1101001111101111;
				18'b000110000100101111: oled_data = 16'b1011001001001001;
				18'b000110000110101111: oled_data = 16'b1011001001001001;
				18'b000110001000101111: oled_data = 16'b1011001001101001;
				18'b000110001010101111: oled_data = 16'b1011001001001001;
				18'b000110001100101111: oled_data = 16'b1011001000101001;
				18'b000110001110101111: oled_data = 16'b1011001000101001;
				18'b000110010000101111: oled_data = 16'b1001100111001000;
				18'b000110010010101111: oled_data = 16'b1000000101000110;
				18'b000110010100101111: oled_data = 16'b1000000100100110;
				18'b000110010110101111: oled_data = 16'b1000000100100101;
				18'b000110011000101111: oled_data = 16'b1001100111000111;
				18'b000110011010101111: oled_data = 16'b1010101000101001;
				18'b000110011100101111: oled_data = 16'b1010001000001000;
				18'b000110011110101111: oled_data = 16'b1001100111100111;
				18'b000110100000101111: oled_data = 16'b1010000111101000;
				18'b000110100010101111: oled_data = 16'b1010100111101000;
				18'b000110100100101111: oled_data = 16'b1010101000001000;
				18'b000110100110101111: oled_data = 16'b1010000111100111;
				18'b000100011000110000: oled_data = 16'b1010101110110001;
				18'b000100011010110000: oled_data = 16'b1100110001010011;
				18'b000100011100110000: oled_data = 16'b1101010010010101;
				18'b000100011110110000: oled_data = 16'b1101010010010101;
				18'b000100100000110000: oled_data = 16'b1101010010010100;
				18'b000100100010110000: oled_data = 16'b1101010010010100;
				18'b000100100100110000: oled_data = 16'b1101110010010100;
				18'b000100100110110000: oled_data = 16'b1101110010010100;
				18'b000100101000110000: oled_data = 16'b1101110010010101;
				18'b000100101010110000: oled_data = 16'b1100110000110011;
				18'b000100101100110000: oled_data = 16'b1010101100101111;
				18'b000100101110110000: oled_data = 16'b1011001101010000;
				18'b000100110000110000: oled_data = 16'b1011001101010000;
				18'b000100110010110000: oled_data = 16'b1010101100110000;
				18'b000100110100110000: oled_data = 16'b1101010001110100;
				18'b000100110110110000: oled_data = 16'b1101110010110101;
				18'b000100111000110000: oled_data = 16'b1101110010010101;
				18'b000100111010110000: oled_data = 16'b1101110010010101;
				18'b000100111100110000: oled_data = 16'b1101110010010101;
				18'b000100111110110000: oled_data = 16'b1101110010010101;
				18'b000101000000110000: oled_data = 16'b1101110010110101;
				18'b000101000010110000: oled_data = 16'b1101110010110101;
				18'b000101000100110000: oled_data = 16'b1101010010010101;
				18'b000101000110110000: oled_data = 16'b1101110111011000;
				18'b000101001000110000: oled_data = 16'b1110111100011011;
				18'b000101001010110000: oled_data = 16'b1110111100011010;
				18'b000101001100110000: oled_data = 16'b1110011100011010;
				18'b000101001110110000: oled_data = 16'b1110011011011001;
				18'b000101010000110000: oled_data = 16'b1101111011011001;
				18'b000101010010110000: oled_data = 16'b1110011011011001;
				18'b000101010100110000: oled_data = 16'b1110011011111010;
				18'b000101010110110000: oled_data = 16'b1110011011011001;
				18'b000101011000110000: oled_data = 16'b1101111010111001;
				18'b000101011010110000: oled_data = 16'b1100110111110110;
				18'b000101011100110000: oled_data = 16'b1100010101110101;
				18'b000101011110110000: oled_data = 16'b1011110011010010;
				18'b000101100000110000: oled_data = 16'b1011010000010000;
				18'b000101100010110000: oled_data = 16'b1011001101101111;
				18'b000101100100110000: oled_data = 16'b1011101110001111;
				18'b000101100110110000: oled_data = 16'b1011101111010000;
				18'b000101101000110000: oled_data = 16'b1011001111010000;
				18'b000101101010110000: oled_data = 16'b1100110001110010;
				18'b000101101100110000: oled_data = 16'b1101110100110101;
				18'b000101101110110000: oled_data = 16'b1101110100110101;
				18'b000101110000110000: oled_data = 16'b1101110100110101;
				18'b000101110010110000: oled_data = 16'b1101010101110101;
				18'b000101110100110000: oled_data = 16'b1110011011011010;
				18'b000101110110110000: oled_data = 16'b1110011011111010;
				18'b000101111000110000: oled_data = 16'b1110011011111010;
				18'b000101111010110000: oled_data = 16'b1110011011111010;
				18'b000101111100110000: oled_data = 16'b1110011100011010;
				18'b000101111110110000: oled_data = 16'b1011101110101110;
				18'b000110000000110000: oled_data = 16'b1011001001101010;
				18'b000110000010110000: oled_data = 16'b1100101110101110;
				18'b000110000100110000: oled_data = 16'b1011001000101001;
				18'b000110000110110000: oled_data = 16'b1011001000101001;
				18'b000110001000110000: oled_data = 16'b1100101101101101;
				18'b000110001010110000: oled_data = 16'b1011101001101010;
				18'b000110001100110000: oled_data = 16'b1011001000101001;
				18'b000110001110110000: oled_data = 16'b1011001001001001;
				18'b000110010000110000: oled_data = 16'b1001100111000111;
				18'b000110010010110000: oled_data = 16'b1000100110100111;
				18'b000110010100110000: oled_data = 16'b1001100111000111;
				18'b000110010110110000: oled_data = 16'b1000000101000101;
				18'b000110011000110000: oled_data = 16'b1000000100100101;
				18'b000110011010110000: oled_data = 16'b1001000110000110;
				18'b000110011100110000: oled_data = 16'b1010000111101000;
				18'b000110011110110000: oled_data = 16'b1010001000001000;
				18'b000110100000110000: oled_data = 16'b1010000111101000;
				18'b000110100010110000: oled_data = 16'b1001100111000111;
				18'b000110100100110000: oled_data = 16'b1001100111000111;
				18'b000110100110110000: oled_data = 16'b1001100111000111;
				18'b000100011000110001: oled_data = 16'b1100110000110011;
				18'b000100011010110001: oled_data = 16'b1101010001110100;
				18'b000100011100110001: oled_data = 16'b1101010001110100;
				18'b000100011110110001: oled_data = 16'b1101010001010100;
				18'b000100100000110001: oled_data = 16'b1101010001110100;
				18'b000100100010110001: oled_data = 16'b1101010001110100;
				18'b000100100100110001: oled_data = 16'b1101010001110100;
				18'b000100100110110001: oled_data = 16'b1101010001110100;
				18'b000100101000110001: oled_data = 16'b1101010010010100;
				18'b000100101010110001: oled_data = 16'b1011101110010001;
				18'b000100101100110001: oled_data = 16'b1010101100001111;
				18'b000100101110110001: oled_data = 16'b1010101100110000;
				18'b000100110000110001: oled_data = 16'b1010101100110000;
				18'b000100110010110001: oled_data = 16'b1011001101110001;
				18'b000100110100110001: oled_data = 16'b1101010001110100;
				18'b000100110110110001: oled_data = 16'b1101110010010100;
				18'b000100111000110001: oled_data = 16'b1101010001110100;
				18'b000100111010110001: oled_data = 16'b1101010001110100;
				18'b000100111100110001: oled_data = 16'b1101010001110100;
				18'b000100111110110001: oled_data = 16'b1101010001110100;
				18'b000101000000110001: oled_data = 16'b1101010010010100;
				18'b000101000010110001: oled_data = 16'b1101010010010100;
				18'b000101000100110001: oled_data = 16'b1101010001110100;
				18'b000101000110110001: oled_data = 16'b1100110101010101;
				18'b000101001000110001: oled_data = 16'b1101110111110111;
				18'b000101001010110001: oled_data = 16'b1101010110110110;
				18'b000101001100110001: oled_data = 16'b1100110111110110;
				18'b000101001110110001: oled_data = 16'b1110011011011001;
				18'b000101010000110001: oled_data = 16'b1110011011011001;
				18'b000101010010110001: oled_data = 16'b1110011011111010;
				18'b000101010100110001: oled_data = 16'b1110011011111010;
				18'b000101010110110001: oled_data = 16'b1110011011111010;
				18'b000101011000110001: oled_data = 16'b1101111010111001;
				18'b000101011010110001: oled_data = 16'b1100110110110101;
				18'b000101011100110001: oled_data = 16'b1011001111110000;
				18'b000101011110110001: oled_data = 16'b1011101110110000;
				18'b000101100000110001: oled_data = 16'b1100001111010000;
				18'b000101100010110001: oled_data = 16'b1011001110001111;
				18'b000101100100110001: oled_data = 16'b1011101110110000;
				18'b000101100110110001: oled_data = 16'b1011101111010000;
				18'b000101101000110001: oled_data = 16'b1100010000110001;
				18'b000101101010110001: oled_data = 16'b1101110100110101;
				18'b000101101100110001: oled_data = 16'b1101110100010101;
				18'b000101101110110001: oled_data = 16'b1101110100110101;
				18'b000101110000110001: oled_data = 16'b1101010100010101;
				18'b000101110010110001: oled_data = 16'b1101010101110110;
				18'b000101110100110001: oled_data = 16'b1110011011111010;
				18'b000101110110110001: oled_data = 16'b1110011011111010;
				18'b000101111000110001: oled_data = 16'b1110011011111010;
				18'b000101111010110001: oled_data = 16'b1110011011011010;
				18'b000101111100110001: oled_data = 16'b1110011100011010;
				18'b000101111110110001: oled_data = 16'b1011101111101111;
				18'b000110000000110001: oled_data = 16'b1011001001001010;
				18'b000110000010110001: oled_data = 16'b1100001101101101;
				18'b000110000100110001: oled_data = 16'b1011001000101001;
				18'b000110000110110001: oled_data = 16'b1011001001001001;
				18'b000110001000110001: oled_data = 16'b1100101101101101;
				18'b000110001010110001: oled_data = 16'b1011001001001001;
				18'b000110001100110001: oled_data = 16'b1011001000101001;
				18'b000110001110110001: oled_data = 16'b1011001000101001;
				18'b000110010000110001: oled_data = 16'b1001000110100111;
				18'b000110010010110001: oled_data = 16'b1001100111000111;
				18'b000110010100110001: oled_data = 16'b1010101000101001;
				18'b000110010110110001: oled_data = 16'b1010000111101000;
				18'b000110011000110001: oled_data = 16'b1001000110000111;
				18'b000110011010110001: oled_data = 16'b1000000100100101;
				18'b000110011100110001: oled_data = 16'b1000000101000101;
				18'b000110011110110001: oled_data = 16'b1001000110000110;
				18'b000110100000110001: oled_data = 16'b1010000111000111;
				18'b000110100010110001: oled_data = 16'b1010000111101000;
				18'b000110100100110001: oled_data = 16'b1010000111001000;
				18'b000110100110110001: oled_data = 16'b1010000111001000;
				18'b000100011000110010: oled_data = 16'b1100110001010011;
				18'b000100011010110010: oled_data = 16'b1101010001010011;
				18'b000100011100110010: oled_data = 16'b1101010001010011;
				18'b000100011110110010: oled_data = 16'b1101010000110011;
				18'b000100100000110010: oled_data = 16'b1101010001010100;
				18'b000100100010110010: oled_data = 16'b1101010001010100;
				18'b000100100100110010: oled_data = 16'b1101010001010100;
				18'b000100100110110010: oled_data = 16'b1100110000110011;
				18'b000100101000110010: oled_data = 16'b1101010001010100;
				18'b000100101010110010: oled_data = 16'b1010101100001111;
				18'b000100101100110010: oled_data = 16'b1010101100001111;
				18'b000100101110110010: oled_data = 16'b1010101100001111;
				18'b000100110000110010: oled_data = 16'b1010101100001111;
				18'b000100110010110010: oled_data = 16'b1100001111110010;
				18'b000100110100110010: oled_data = 16'b1101010001010100;
				18'b000100110110110010: oled_data = 16'b1101010001110100;
				18'b000100111000110010: oled_data = 16'b1101010001110100;
				18'b000100111010110010: oled_data = 16'b1101010001110100;
				18'b000100111100110010: oled_data = 16'b1101010001110100;
				18'b000100111110110010: oled_data = 16'b1101010001110100;
				18'b000101000000110010: oled_data = 16'b1101010001110100;
				18'b000101000010110010: oled_data = 16'b1101010001110100;
				18'b000101000100110010: oled_data = 16'b1100110001010011;
				18'b000101000110110010: oled_data = 16'b1100010000110010;
				18'b000101001000110010: oled_data = 16'b1011110000110010;
				18'b000101001010110010: oled_data = 16'b1011110001010010;
				18'b000101001100110010: oled_data = 16'b1101111000111000;
				18'b000101001110110010: oled_data = 16'b1110011011011010;
				18'b000101010000110010: oled_data = 16'b1110011011011001;
				18'b000101010010110010: oled_data = 16'b1110011011011001;
				18'b000101010100110010: oled_data = 16'b1110011011011001;
				18'b000101010110110010: oled_data = 16'b1110011011011001;
				18'b000101011000110010: oled_data = 16'b1110011011111010;
				18'b000101011010110010: oled_data = 16'b1110011011011001;
				18'b000101011100110010: oled_data = 16'b1100110100110100;
				18'b000101011110110010: oled_data = 16'b1011001111110000;
				18'b000101100000110010: oled_data = 16'b1011101111010000;
				18'b000101100010110010: oled_data = 16'b1011001110001111;
				18'b000101100100110010: oled_data = 16'b1100001111110001;
				18'b000101100110110010: oled_data = 16'b1100110001010010;
				18'b000101101000110010: oled_data = 16'b1101010011110100;
				18'b000101101010110010: oled_data = 16'b1101110100010101;
				18'b000101101100110010: oled_data = 16'b1101110100010101;
				18'b000101101110110010: oled_data = 16'b1101110100010101;
				18'b000101110000110010: oled_data = 16'b1101010011110100;
				18'b000101110010110010: oled_data = 16'b1101110110010110;
				18'b000101110100110010: oled_data = 16'b1110011011011010;
				18'b000101110110110010: oled_data = 16'b1110011011011010;
				18'b000101111000110010: oled_data = 16'b1110011011011010;
				18'b000101111010110010: oled_data = 16'b1110011011011010;
				18'b000101111100110010: oled_data = 16'b1110011011111010;
				18'b000101111110110010: oled_data = 16'b1011001111001110;
				18'b000110000000110010: oled_data = 16'b1011001001001001;
				18'b000110000010110010: oled_data = 16'b1011101100101101;
				18'b000110000100110010: oled_data = 16'b1011001000101001;
				18'b000110000110110010: oled_data = 16'b1011001001001001;
				18'b000110001000110010: oled_data = 16'b1011101010101011;
				18'b000110001010110010: oled_data = 16'b1011001000101001;
				18'b000110001100110010: oled_data = 16'b1011001000101000;
				18'b000110001110110010: oled_data = 16'b1011001000101001;
				18'b000110010000110010: oled_data = 16'b1001000110100111;
				18'b000110010010110010: oled_data = 16'b1010000111000111;
				18'b000110010100110010: oled_data = 16'b1010101000001000;
				18'b000110010110110010: oled_data = 16'b1010101000001000;
				18'b000110011000110010: oled_data = 16'b1010101000001000;
				18'b000110011010110010: oled_data = 16'b1010000111101000;
				18'b000110011100110010: oled_data = 16'b1010000111001000;
				18'b000110011110110010: oled_data = 16'b1010000111000111;
				18'b000110100000110010: oled_data = 16'b1010000111000111;
				18'b000110100010110010: oled_data = 16'b1010000111000111;
				18'b000110100100110010: oled_data = 16'b1010000111000111;
				18'b000110100110110010: oled_data = 16'b1010000111000111;
				18'b000100011000110011: oled_data = 16'b1100110000010011;
				18'b000100011010110011: oled_data = 16'b1100110000010011;
				18'b000100011100110011: oled_data = 16'b1101010000110011;
				18'b000100011110110011: oled_data = 16'b1100110000010011;
				18'b000100100000110011: oled_data = 16'b1101010000110011;
				18'b000100100010110011: oled_data = 16'b1100110000110011;
				18'b000100100100110011: oled_data = 16'b1100101111110010;
				18'b000100100110110011: oled_data = 16'b1100101111110010;
				18'b000100101000110011: oled_data = 16'b1100001111110010;
				18'b000100101010110011: oled_data = 16'b1010001010101110;
				18'b000100101100110011: oled_data = 16'b1010001011101111;
				18'b000100101110110011: oled_data = 16'b1010001011101111;
				18'b000100110000110011: oled_data = 16'b1011001101010000;
				18'b000100110010110011: oled_data = 16'b1100010000010011;
				18'b000100110100110011: oled_data = 16'b1101010001010100;
				18'b000100110110110011: oled_data = 16'b1101010001010100;
				18'b000100111000110011: oled_data = 16'b1101010001010011;
				18'b000100111010110011: oled_data = 16'b1101010001010011;
				18'b000100111100110011: oled_data = 16'b1101010001010100;
				18'b000100111110110011: oled_data = 16'b1101010001010100;
				18'b000101000000110011: oled_data = 16'b1101010001010100;
				18'b000101000010110011: oled_data = 16'b1101010001010100;
				18'b000101000100110011: oled_data = 16'b1100010000010010;
				18'b000101000110110011: oled_data = 16'b1100010000110010;
				18'b000101001000110011: oled_data = 16'b1100010000110010;
				18'b000101001010110011: oled_data = 16'b1101010101010110;
				18'b000101001100110011: oled_data = 16'b1110011010011001;
				18'b000101001110110011: oled_data = 16'b1110011010111001;
				18'b000101010000110011: oled_data = 16'b1101111010111001;
				18'b000101010010110011: oled_data = 16'b1101111010111001;
				18'b000101010100110011: oled_data = 16'b1101111010111001;
				18'b000101010110110011: oled_data = 16'b1110011010111001;
				18'b000101011000110011: oled_data = 16'b1110011010111001;
				18'b000101011010110011: oled_data = 16'b1110011010111001;
				18'b000101011100110011: oled_data = 16'b1101111000110111;
				18'b000101011110110011: oled_data = 16'b1100010010110010;
				18'b000101100000110011: oled_data = 16'b1100010001010010;
				18'b000101100010110011: oled_data = 16'b1100010001010010;
				18'b000101100100110011: oled_data = 16'b1101010010110011;
				18'b000101100110110011: oled_data = 16'b1101010011010011;
				18'b000101101000110011: oled_data = 16'b1101010011010100;
				18'b000101101010110011: oled_data = 16'b1101010011110100;
				18'b000101101100110011: oled_data = 16'b1101010011110100;
				18'b000101101110110011: oled_data = 16'b1101010011110100;
				18'b000101110000110011: oled_data = 16'b1101010011010100;
				18'b000101110010110011: oled_data = 16'b1101110100110101;
				18'b000101110100110011: oled_data = 16'b1101111000111000;
				18'b000101110110110011: oled_data = 16'b1101111010111001;
				18'b000101111000110011: oled_data = 16'b1110011010111001;
				18'b000101111010110011: oled_data = 16'b1101111010011001;
				18'b000101111100110011: oled_data = 16'b1101111011011001;
				18'b000101111110110011: oled_data = 16'b1011001111001110;
				18'b000110000000110011: oled_data = 16'b1011001001001001;
				18'b000110000010110011: oled_data = 16'b1011101100001100;
				18'b000110000100110011: oled_data = 16'b1011001000001001;
				18'b000110000110110011: oled_data = 16'b1011001000101001;
				18'b000110001000110011: oled_data = 16'b1011001000001000;
				18'b000110001010110011: oled_data = 16'b1011001000001000;
				18'b000110001100110011: oled_data = 16'b1010101000001000;
				18'b000110001110110011: oled_data = 16'b1010101000001000;
				18'b000110010000110011: oled_data = 16'b1000100110000110;
				18'b000110010010110011: oled_data = 16'b1010000111101000;
				18'b000110010100110011: oled_data = 16'b1010100111101000;
				18'b000110010110110011: oled_data = 16'b1010100111101000;
				18'b000110011000110011: oled_data = 16'b1010000111101000;
				18'b000110011010110011: oled_data = 16'b1010000111101000;
				18'b000110011100110011: oled_data = 16'b1010000111000111;
				18'b000110011110110011: oled_data = 16'b1010000111000111;
				18'b000110100000110011: oled_data = 16'b1010000111000111;
				18'b000110100010110011: oled_data = 16'b1001100111000111;
				18'b000110100100110011: oled_data = 16'b1001100111000111;
				18'b000110100110110011: oled_data = 16'b1001100111000111;
				18'b000100011000110100: oled_data = 16'b1100101111110010;
				18'b000100011010110100: oled_data = 16'b1100101111110011;
				18'b000100011100110100: oled_data = 16'b1100101111110010;
				18'b000100011110110100: oled_data = 16'b1100110000010010;
				18'b000100100000110100: oled_data = 16'b1100110000010011;
				18'b000100100010110100: oled_data = 16'b1100101111110010;
				18'b000100100100110100: oled_data = 16'b1011101101110000;
				18'b000100100110110100: oled_data = 16'b1100110000010010;
				18'b000100101000110100: oled_data = 16'b1011001101001111;
				18'b000100101010110100: oled_data = 16'b1001101010101110;
				18'b000100101100110100: oled_data = 16'b1010001011101110;
				18'b000100101110110100: oled_data = 16'b1001101011001110;
				18'b000100110000110100: oled_data = 16'b1011101110010001;
				18'b000100110010110100: oled_data = 16'b1100001111110010;
				18'b000100110100110100: oled_data = 16'b1100110000110011;
				18'b000100110110110100: oled_data = 16'b1101010000110011;
				18'b000100111000110100: oled_data = 16'b1100110000110011;
				18'b000100111010110100: oled_data = 16'b1100110000110011;
				18'b000100111100110100: oled_data = 16'b1100110000110011;
				18'b000100111110110100: oled_data = 16'b1100110000110011;
				18'b000101000000110100: oled_data = 16'b1100110000110011;
				18'b000101000010110100: oled_data = 16'b1100110000110011;
				18'b000101000100110100: oled_data = 16'b1100001111110001;
				18'b000101000110110100: oled_data = 16'b1100010000110010;
				18'b000101001000110100: oled_data = 16'b1100010001010010;
				18'b000101001010110100: oled_data = 16'b1100110100010100;
				18'b000101001100110100: oled_data = 16'b1101011001011000;
				18'b000101001110110100: oled_data = 16'b1101111010011001;
				18'b000101010000110100: oled_data = 16'b1101111010011001;
				18'b000101010010110100: oled_data = 16'b1110011010111001;
				18'b000101010100110100: oled_data = 16'b1110011010111001;
				18'b000101010110110100: oled_data = 16'b1110011010111001;
				18'b000101011000110100: oled_data = 16'b1110011010111001;
				18'b000101011010110100: oled_data = 16'b1101111010111001;
				18'b000101011100110100: oled_data = 16'b1101111001111000;
				18'b000101011110110100: oled_data = 16'b1100110101010100;
				18'b000101100000110100: oled_data = 16'b1100110010110011;
				18'b000101100010110100: oled_data = 16'b1100110001110010;
				18'b000101100100110100: oled_data = 16'b1101010011010011;
				18'b000101100110110100: oled_data = 16'b1101010011010011;
				18'b000101101000110100: oled_data = 16'b1101010011010100;
				18'b000101101010110100: oled_data = 16'b1101010011010100;
				18'b000101101100110100: oled_data = 16'b1101010011010100;
				18'b000101101110110100: oled_data = 16'b1101010011010100;
				18'b000101110000110100: oled_data = 16'b1101010011010100;
				18'b000101110010110100: oled_data = 16'b1100010010010010;
				18'b000101110100110100: oled_data = 16'b1001110000010000;
				18'b000101110110110100: oled_data = 16'b1100111000010111;
				18'b000101111000110100: oled_data = 16'b1101011000110111;
				18'b000101111010110100: oled_data = 16'b1100010111110110;
				18'b000101111100110100: oled_data = 16'b1101011001010111;
				18'b000101111110110100: oled_data = 16'b1011001110001101;
				18'b000110000000110100: oled_data = 16'b1011001000101001;
				18'b000110000010110100: oled_data = 16'b1011001011001011;
				18'b000110000100110100: oled_data = 16'b1011001000001000;
				18'b000110000110110100: oled_data = 16'b1011001000001000;
				18'b000110001000110100: oled_data = 16'b1010101000001000;
				18'b000110001010110100: oled_data = 16'b1010101000001000;
				18'b000110001100110100: oled_data = 16'b1010101000001000;
				18'b000110001110110100: oled_data = 16'b1010101000001000;
				18'b000110010000110100: oled_data = 16'b1000100101100110;
				18'b000110010010110100: oled_data = 16'b1010000111101000;
				18'b000110010100110100: oled_data = 16'b1010100111101000;
				18'b000110010110110100: oled_data = 16'b1010000111100111;
				18'b000110011000110100: oled_data = 16'b1010000111100111;
				18'b000110011010110100: oled_data = 16'b1010000111000111;
				18'b000110011100110100: oled_data = 16'b1010000111000111;
				18'b000110011110110100: oled_data = 16'b1010000111000111;
				18'b000110100000110100: oled_data = 16'b1001100111000111;
				18'b000110100010110100: oled_data = 16'b1001100111000111;
				18'b000110100100110100: oled_data = 16'b1001100111000111;
				18'b000110100110110100: oled_data = 16'b1001100110100110;
				18'b000100011000110101: oled_data = 16'b1100001111010010;
				18'b000100011010110101: oled_data = 16'b1100001111010010;
				18'b000100011100110101: oled_data = 16'b1100001111110001;
				18'b000100011110110101: oled_data = 16'b1100001111110010;
				18'b000100100000110101: oled_data = 16'b1100101111110010;
				18'b000100100010110101: oled_data = 16'b1011001101010000;
				18'b000100100100110101: oled_data = 16'b1011101101110000;
				18'b000100100110110101: oled_data = 16'b1100001111110010;
				18'b000100101000110101: oled_data = 16'b1001101010101101;
				18'b000100101010110101: oled_data = 16'b1001101010101110;
				18'b000100101100110101: oled_data = 16'b1001101011001110;
				18'b000100101110110101: oled_data = 16'b1010001011001110;
				18'b000100110000110101: oled_data = 16'b1100001111010010;
				18'b000100110010110101: oled_data = 16'b1100001110110001;
				18'b000100110100110101: oled_data = 16'b1100110000010011;
				18'b000100110110110101: oled_data = 16'b1100110000010011;
				18'b000100111000110101: oled_data = 16'b1100110000010011;
				18'b000100111010110101: oled_data = 16'b1100110000010011;
				18'b000100111100110101: oled_data = 16'b1100101111110011;
				18'b000100111110110101: oled_data = 16'b1100101111110011;
				18'b000101000000110101: oled_data = 16'b1100110000010011;
				18'b000101000010110101: oled_data = 16'b1100110000010010;
				18'b000101000100110101: oled_data = 16'b1011110000010010;
				18'b000101000110110101: oled_data = 16'b1100010000110010;
				18'b000101001000110101: oled_data = 16'b1100010001110011;
				18'b000101001010110101: oled_data = 16'b1100110100110100;
				18'b000101001100110101: oled_data = 16'b1101011001011000;
				18'b000101001110110101: oled_data = 16'b1101111010011000;
				18'b000101010000110101: oled_data = 16'b1101111010011000;
				18'b000101010010110101: oled_data = 16'b1101111001111000;
				18'b000101010100110101: oled_data = 16'b1101111010011000;
				18'b000101010110110101: oled_data = 16'b1101111010011000;
				18'b000101011000110101: oled_data = 16'b1101111010011000;
				18'b000101011010110101: oled_data = 16'b1101111010011001;
				18'b000101011100110101: oled_data = 16'b1101111001111000;
				18'b000101011110110101: oled_data = 16'b1100110101010101;
				18'b000101100000110101: oled_data = 16'b1100110010010011;
				18'b000101100010110101: oled_data = 16'b1100010000110001;
				18'b000101100100110101: oled_data = 16'b1101010010110011;
				18'b000101100110110101: oled_data = 16'b1101010010110011;
				18'b000101101000110101: oled_data = 16'b1101010010010100;
				18'b000101101010110101: oled_data = 16'b1100110010110011;
				18'b000101101100110101: oled_data = 16'b1100110010110011;
				18'b000101101110110101: oled_data = 16'b1101010010010100;
				18'b000101110000110101: oled_data = 16'b1101010010110100;
				18'b000101110010110101: oled_data = 16'b1010001111001111;
				18'b000101110100110101: oled_data = 16'b0010100011100011;
				18'b000101110110110101: oled_data = 16'b0110101100001011;
				18'b000101111000110101: oled_data = 16'b1010010010110001;
				18'b000101111010110101: oled_data = 16'b1010010011010010;
				18'b000101111100110101: oled_data = 16'b1011010100010011;
				18'b000101111110110101: oled_data = 16'b1010001100001100;
				18'b000110000000110101: oled_data = 16'b1010101000001000;
				18'b000110000010110101: oled_data = 16'b1011001010001010;
				18'b000110000100110101: oled_data = 16'b1010100111101000;
				18'b000110000110110101: oled_data = 16'b1010101000001000;
				18'b000110001000110101: oled_data = 16'b1010100111101000;
				18'b000110001010110101: oled_data = 16'b1010100111101000;
				18'b000110001100110101: oled_data = 16'b1010100111101000;
				18'b000110001110110101: oled_data = 16'b1010000111101000;
				18'b000110010000110101: oled_data = 16'b1000100101100110;
				18'b000110010010110101: oled_data = 16'b1010000111001000;
				18'b000110010100110101: oled_data = 16'b1010000111001000;
				18'b000110010110110101: oled_data = 16'b1010000111000111;
				18'b000110011000110101: oled_data = 16'b1001100111000111;
				18'b000110011010110101: oled_data = 16'b1010000111000111;
				18'b000110011100110101: oled_data = 16'b1001100111000111;
				18'b000110011110110101: oled_data = 16'b1001100111000111;
				18'b000110100000110101: oled_data = 16'b1001100110100111;
				18'b000110100010110101: oled_data = 16'b1001100110100110;
				18'b000110100100110101: oled_data = 16'b1001100110100111;
				18'b000110100110110101: oled_data = 16'b1001100110100111;
				18'b000100011000110110: oled_data = 16'b1100001110110010;
				18'b000100011010110110: oled_data = 16'b1100001110110010;
				18'b000100011100110110: oled_data = 16'b1100001111010001;
				18'b000100011110110110: oled_data = 16'b1100001111010001;
				18'b000100100000110110: oled_data = 16'b1011101110010001;
				18'b000100100010110110: oled_data = 16'b1010001011001110;
				18'b000100100100110110: oled_data = 16'b1100001110110010;
				18'b000100100110110110: oled_data = 16'b1011001101110000;
				18'b000100101000110110: oled_data = 16'b1001001010001101;
				18'b000100101010110110: oled_data = 16'b1001001010001101;
				18'b000100101100110110: oled_data = 16'b1001101010001101;
				18'b000100101110110110: oled_data = 16'b1001101010101110;
				18'b000100110000110110: oled_data = 16'b1011101110110001;
				18'b000100110010110110: oled_data = 16'b1100001110110001;
				18'b000100110100110110: oled_data = 16'b1100101111110010;
				18'b000100110110110110: oled_data = 16'b1100101111110010;
				18'b000100111000110110: oled_data = 16'b1100101111110010;
				18'b000100111010110110: oled_data = 16'b1100001111110010;
				18'b000100111100110110: oled_data = 16'b1100101111110010;
				18'b000100111110110110: oled_data = 16'b1100101111110010;
				18'b000101000000110110: oled_data = 16'b1100101111110010;
				18'b000101000010110110: oled_data = 16'b1100001111010001;
				18'b000101000100110110: oled_data = 16'b1100010000110010;
				18'b000101000110110110: oled_data = 16'b1100010000110010;
				18'b000101001000110110: oled_data = 16'b1100110001110011;
				18'b000101001010110110: oled_data = 16'b1100110101010101;
				18'b000101001100110110: oled_data = 16'b1101011001011000;
				18'b000101001110110110: oled_data = 16'b1101011001111000;
				18'b000101010000110110: oled_data = 16'b1101011001111000;
				18'b000101010010110110: oled_data = 16'b1101011001111000;
				18'b000101010100110110: oled_data = 16'b1101011001111000;
				18'b000101010110110110: oled_data = 16'b1101011001111000;
				18'b000101011000110110: oled_data = 16'b1101011001111000;
				18'b000101011010110110: oled_data = 16'b1101011001111000;
				18'b000101011100110110: oled_data = 16'b1101011001011000;
				18'b000101011110110110: oled_data = 16'b1100110100110100;
				18'b000101100000110110: oled_data = 16'b1100010001010010;
				18'b000101100010110110: oled_data = 16'b1100010000110001;
				18'b000101100100110110: oled_data = 16'b1100110010010011;
				18'b000101100110110110: oled_data = 16'b1100110010010011;
				18'b000101101000110110: oled_data = 16'b1100110001110011;
				18'b000101101010110110: oled_data = 16'b1100110010010011;
				18'b000101101100110110: oled_data = 16'b1100110010010010;
				18'b000101101110110110: oled_data = 16'b1100110010010011;
				18'b000101110000110110: oled_data = 16'b1101010010010100;
				18'b000101110010110110: oled_data = 16'b0110101000101001;
				18'b000101110100110110: oled_data = 16'b0001100010000001;
				18'b000101110110110110: oled_data = 16'b0010100011000010;
				18'b000101111000110110: oled_data = 16'b0100000101100101;
				18'b000101111010110110: oled_data = 16'b0111001010101010;
				18'b000101111100110110: oled_data = 16'b1001001110001101;
				18'b000101111110110110: oled_data = 16'b1010001010101010;
				18'b000110000000110110: oled_data = 16'b1010100111101000;
				18'b000110000010110110: oled_data = 16'b1010101001001001;
				18'b000110000100110110: oled_data = 16'b1010100111101000;
				18'b000110000110110110: oled_data = 16'b1010100111101000;
				18'b000110001000110110: oled_data = 16'b1010100111100111;
				18'b000110001010110110: oled_data = 16'b1010000111100111;
				18'b000110001100110110: oled_data = 16'b1010100111000111;
				18'b000110001110110110: oled_data = 16'b1001100111000111;
				18'b000110010000110110: oled_data = 16'b1000100101100110;
				18'b000110010010110110: oled_data = 16'b1010000111001000;
				18'b000110010100110110: oled_data = 16'b1010000111000111;
				18'b000110010110110110: oled_data = 16'b1001100111000111;
				18'b000110011000110110: oled_data = 16'b1001100110100111;
				18'b000110011010110110: oled_data = 16'b1001100110100111;
				18'b000110011100110110: oled_data = 16'b1001100110100111;
				18'b000110011110110110: oled_data = 16'b1001100110100111;
				18'b000110100000110110: oled_data = 16'b1001100110100110;
				18'b000110100010110110: oled_data = 16'b1001100110100110;
				18'b000110100100110110: oled_data = 16'b1001000110100110;
				18'b000110100110110110: oled_data = 16'b1001000110000110;
				18'b000100011000110111: oled_data = 16'b1011101110110001;
				18'b000100011010110111: oled_data = 16'b1100001110010001;
				18'b000100011100110111: oled_data = 16'b1100001110010001;
				18'b000100011110110111: oled_data = 16'b1100001110110001;
				18'b000100100000110111: oled_data = 16'b1010001011001110;
				18'b000100100010110111: oled_data = 16'b1010101011101111;
				18'b000100100100110111: oled_data = 16'b1100001110110010;
				18'b000100100110110111: oled_data = 16'b1010001011001110;
				18'b000100101000110111: oled_data = 16'b1001001001101100;
				18'b000100101010110111: oled_data = 16'b1001001010001101;
				18'b000100101100110111: oled_data = 16'b1001001001101101;
				18'b000100101110110111: oled_data = 16'b1001101011001110;
				18'b000100110000110111: oled_data = 16'b1011101110010001;
				18'b000100110010110111: oled_data = 16'b1100001110110001;
				18'b000100110100110111: oled_data = 16'b1100001111010010;
				18'b000100110110110111: oled_data = 16'b1100001111010010;
				18'b000100111000110111: oled_data = 16'b1100001111010010;
				18'b000100111010110111: oled_data = 16'b1100001111010010;
				18'b000100111100110111: oled_data = 16'b1100001111010010;
				18'b000100111110110111: oled_data = 16'b1100001111010010;
				18'b000101000000110111: oled_data = 16'b1100001111010010;
				18'b000101000010110111: oled_data = 16'b1011101110110001;
				18'b000101000100110111: oled_data = 16'b1100010000110010;
				18'b000101000110110111: oled_data = 16'b1100110001110011;
				18'b000101001000110111: oled_data = 16'b1100010001110010;
				18'b000101001010110111: oled_data = 16'b1100110101010101;
				18'b000101001100110111: oled_data = 16'b1101011001010111;
				18'b000101001110110111: oled_data = 16'b1101011001010111;
				18'b000101010000110111: oled_data = 16'b1101011001010111;
				18'b000101010010110111: oled_data = 16'b1101011001010111;
				18'b000101010100110111: oled_data = 16'b1101011001010111;
				18'b000101010110110111: oled_data = 16'b1101011001011000;
				18'b000101011000110111: oled_data = 16'b1101011001011000;
				18'b000101011010110111: oled_data = 16'b1101011001011000;
				18'b000101011100110111: oled_data = 16'b1101011000110111;
				18'b000101011110110111: oled_data = 16'b1100010100010100;
				18'b000101100000110111: oled_data = 16'b1100010001010001;
				18'b000101100010110111: oled_data = 16'b1100010000010001;
				18'b000101100100110111: oled_data = 16'b1100110001110010;
				18'b000101100110110111: oled_data = 16'b1100110001110010;
				18'b000101101000110111: oled_data = 16'b1100110001110010;
				18'b000101101010110111: oled_data = 16'b1100110001110010;
				18'b000101101100110111: oled_data = 16'b1100110001110010;
				18'b000101101110110111: oled_data = 16'b1100110001110010;
				18'b000101110000110111: oled_data = 16'b1011101111110001;
				18'b000101110010110111: oled_data = 16'b0011100100000100;
				18'b000101110100110111: oled_data = 16'b0011000011100011;
				18'b000101110110110111: oled_data = 16'b0101000110000101;
				18'b000101111000110111: oled_data = 16'b0111001001000110;
				18'b000101111010110111: oled_data = 16'b0111101010000111;
				18'b000101111100110111: oled_data = 16'b0111101001100110;
				18'b000101111110110111: oled_data = 16'b1000101000100111;
				18'b000110000000110111: oled_data = 16'b1010100111101000;
				18'b000110000010110111: oled_data = 16'b1010101000101000;
				18'b000110000100110111: oled_data = 16'b1010100111101000;
				18'b000110000110110111: oled_data = 16'b1010100111100111;
				18'b000110001000110111: oled_data = 16'b1010000111100111;
				18'b000110001010110111: oled_data = 16'b1010000111100111;
				18'b000110001100110111: oled_data = 16'b1010000111000111;
				18'b000110001110110111: oled_data = 16'b1001100110100110;
				18'b000110010000110111: oled_data = 16'b1000100110000110;
				18'b000110010010110111: oled_data = 16'b1010000110100111;
				18'b000110010100110111: oled_data = 16'b1010000110100111;
				18'b000110010110110111: oled_data = 16'b1001100110100111;
				18'b000110011000110111: oled_data = 16'b1001000110100111;
				18'b000110011010110111: oled_data = 16'b1001100110100111;
				18'b000110011100110111: oled_data = 16'b1001100110100111;
				18'b000110011110110111: oled_data = 16'b1001000110100110;
				18'b000110100000110111: oled_data = 16'b1001000110100110;
				18'b000110100010110111: oled_data = 16'b1001000110100110;
				18'b000110100100110111: oled_data = 16'b1001000110000110;
				18'b000110100110110111: oled_data = 16'b1001000110000110;
				18'b001000011000001000: oled_data = 16'b1001101111101011;
				18'b001000011010001000: oled_data = 16'b1010010000001011;
				18'b001000011100001000: oled_data = 16'b1010010000101011;
				18'b001000011110001000: oled_data = 16'b1010110001001011;
				18'b001000100000001000: oled_data = 16'b1010010000101011;
				18'b001000100010001000: oled_data = 16'b1101010111110110;
				18'b001000100100001000: oled_data = 16'b1111011010111011;
				18'b001000100110001000: oled_data = 16'b1110010100110111;
				18'b001000101000001000: oled_data = 16'b1101110011010101;
				18'b001000101010001000: oled_data = 16'b1110010011010110;
				18'b001000101100001000: oled_data = 16'b1101110011010101;
				18'b001000101110001000: oled_data = 16'b1101110011010101;
				18'b001000110000001000: oled_data = 16'b1101110011010101;
				18'b001000110010001000: oled_data = 16'b1101110011010101;
				18'b001000110100001000: oled_data = 16'b1101110011010101;
				18'b001000110110001000: oled_data = 16'b1101110011010101;
				18'b001000111000001000: oled_data = 16'b1101110011010101;
				18'b001000111010001000: oled_data = 16'b1101110011010101;
				18'b001000111100001000: oled_data = 16'b1101110011010101;
				18'b001000111110001000: oled_data = 16'b1101110011010101;
				18'b001001000000001000: oled_data = 16'b1101110011010101;
				18'b001001000010001000: oled_data = 16'b1101110011010101;
				18'b001001000100001000: oled_data = 16'b1101110011010101;
				18'b001001000110001000: oled_data = 16'b1101110011010101;
				18'b001001001000001000: oled_data = 16'b1101110011010101;
				18'b001001001010001000: oled_data = 16'b1101110011010101;
				18'b001001001100001000: oled_data = 16'b1101110011010101;
				18'b001001001110001000: oled_data = 16'b1101110011010101;
				18'b001001010000001000: oled_data = 16'b1101110011010101;
				18'b001001010010001000: oled_data = 16'b1101110011010101;
				18'b001001010100001000: oled_data = 16'b1101110011010101;
				18'b001001010110001000: oled_data = 16'b1101110011010101;
				18'b001001011000001000: oled_data = 16'b1101110011010101;
				18'b001001011010001000: oled_data = 16'b1101110011010101;
				18'b001001011100001000: oled_data = 16'b1101110011010101;
				18'b001001011110001000: oled_data = 16'b1101110011010101;
				18'b001001100000001000: oled_data = 16'b1101110011010101;
				18'b001001100010001000: oled_data = 16'b1101110011010101;
				18'b001001100100001000: oled_data = 16'b1101110011010101;
				18'b001001100110001000: oled_data = 16'b1101110011010101;
				18'b001001101000001000: oled_data = 16'b1101110011010101;
				18'b001001101010001000: oled_data = 16'b1101110011010101;
				18'b001001101100001000: oled_data = 16'b1101110011010101;
				18'b001001101110001000: oled_data = 16'b1101110011010110;
				18'b001001110000001000: oled_data = 16'b1101110010110101;
				18'b001001110010001000: oled_data = 16'b1101010010010100;
				18'b001001110100001000: oled_data = 16'b1110010011110110;
				18'b001001110110001000: oled_data = 16'b1101110011110110;
				18'b001001111000001000: oled_data = 16'b1110010011110110;
				18'b001001111010001000: oled_data = 16'b1101010010010101;
				18'b001001111100001000: oled_data = 16'b1101010010010101;
				18'b001001111110001000: oled_data = 16'b1101110011010110;
				18'b001010000000001000: oled_data = 16'b1101110011010101;
				18'b001010000010001000: oled_data = 16'b1101010010010101;
				18'b001010000100001000: oled_data = 16'b1110011000011001;
				18'b001010000110001000: oled_data = 16'b1101011000011000;
				18'b001010001000001000: oled_data = 16'b0101101001000111;
				18'b001010001010001000: oled_data = 16'b0101101001000110;
				18'b001010001100001000: oled_data = 16'b0111001011000110;
				18'b001010001110001000: oled_data = 16'b0111101100000111;
				18'b001010010000001000: oled_data = 16'b0111101100000111;
				18'b001010010010001000: oled_data = 16'b0111101100000111;
				18'b001010010100001000: oled_data = 16'b0111001100001000;
				18'b001010010110001000: oled_data = 16'b0111001011101000;
				18'b001010011000001000: oled_data = 16'b0110101011101000;
				18'b001010011010001000: oled_data = 16'b0110001011001000;
				18'b001010011100001000: oled_data = 16'b0110001010101000;
				18'b001010011110001000: oled_data = 16'b0101101010001000;
				18'b001010100000001000: oled_data = 16'b0101101010001000;
				18'b001010100010001000: oled_data = 16'b0101001001101000;
				18'b001010100100001000: oled_data = 16'b0101001001001000;
				18'b001010100110001000: oled_data = 16'b0101001001101000;
				18'b001000011000001001: oled_data = 16'b1011010001101011;
				18'b001000011010001001: oled_data = 16'b1011010001101011;
				18'b001000011100001001: oled_data = 16'b1011010001001011;
				18'b001000011110001001: oled_data = 16'b1010110000101011;
				18'b001000100000001001: oled_data = 16'b1011010010101110;
				18'b001000100010001001: oled_data = 16'b1111011010111011;
				18'b001000100100001001: oled_data = 16'b1110010111011001;
				18'b001000100110001001: oled_data = 16'b1101110011010110;
				18'b001000101000001001: oled_data = 16'b1101110011010101;
				18'b001000101010001001: oled_data = 16'b1101110011010101;
				18'b001000101100001001: oled_data = 16'b1101110011010101;
				18'b001000101110001001: oled_data = 16'b1101110011010101;
				18'b001000110000001001: oled_data = 16'b1101110011010101;
				18'b001000110010001001: oled_data = 16'b1101110011010101;
				18'b001000110100001001: oled_data = 16'b1101110011010101;
				18'b001000110110001001: oled_data = 16'b1101110011010101;
				18'b001000111000001001: oled_data = 16'b1101110011010101;
				18'b001000111010001001: oled_data = 16'b1101110011010101;
				18'b001000111100001001: oled_data = 16'b1101110011010101;
				18'b001000111110001001: oled_data = 16'b1101110011010101;
				18'b001001000000001001: oled_data = 16'b1101110011010101;
				18'b001001000010001001: oled_data = 16'b1101110011010101;
				18'b001001000100001001: oled_data = 16'b1101110011010101;
				18'b001001000110001001: oled_data = 16'b1101110011010101;
				18'b001001001000001001: oled_data = 16'b1101110011010101;
				18'b001001001010001001: oled_data = 16'b1101110011010101;
				18'b001001001100001001: oled_data = 16'b1101110011010101;
				18'b001001001110001001: oled_data = 16'b1101110011010101;
				18'b001001010000001001: oled_data = 16'b1101110011010101;
				18'b001001010010001001: oled_data = 16'b1101110011010101;
				18'b001001010100001001: oled_data = 16'b1101110011010101;
				18'b001001010110001001: oled_data = 16'b1101110011010110;
				18'b001001011000001001: oled_data = 16'b1101110010110101;
				18'b001001011010001001: oled_data = 16'b1101110010110101;
				18'b001001011100001001: oled_data = 16'b1101110011010101;
				18'b001001011110001001: oled_data = 16'b1101110011010101;
				18'b001001100000001001: oled_data = 16'b1101110011010101;
				18'b001001100010001001: oled_data = 16'b1101110011010101;
				18'b001001100100001001: oled_data = 16'b1101110011010101;
				18'b001001100110001001: oled_data = 16'b1101110011010101;
				18'b001001101000001001: oled_data = 16'b1101110011010101;
				18'b001001101010001001: oled_data = 16'b1101010001110100;
				18'b001001101100001001: oled_data = 16'b1101110011010101;
				18'b001001101110001001: oled_data = 16'b1101110011010101;
				18'b001001110000001001: oled_data = 16'b1101110011010110;
				18'b001001110010001001: oled_data = 16'b1101010001110100;
				18'b001001110100001001: oled_data = 16'b1101110011010110;
				18'b001001110110001001: oled_data = 16'b1101110011110110;
				18'b001001111000001001: oled_data = 16'b1101110011110110;
				18'b001001111010001001: oled_data = 16'b1101110011010101;
				18'b001001111100001001: oled_data = 16'b1101010001110100;
				18'b001001111110001001: oled_data = 16'b1101110011010110;
				18'b001010000000001001: oled_data = 16'b1101110011010101;
				18'b001010000010001001: oled_data = 16'b1101110010110101;
				18'b001010000100001001: oled_data = 16'b1101110101010111;
				18'b001010000110001001: oled_data = 16'b1111011011111100;
				18'b001010001000001001: oled_data = 16'b1000101110001101;
				18'b001010001010001001: oled_data = 16'b0101101000000101;
				18'b001010001100001001: oled_data = 16'b0111001011000111;
				18'b001010001110001001: oled_data = 16'b0111101100000111;
				18'b001010010000001001: oled_data = 16'b0111101100100111;
				18'b001010010010001001: oled_data = 16'b1000001100101000;
				18'b001010010100001001: oled_data = 16'b1000001100101000;
				18'b001010010110001001: oled_data = 16'b1000101101001000;
				18'b001010011000001001: oled_data = 16'b1000101101101000;
				18'b001010011010001001: oled_data = 16'b1000101101101000;
				18'b001010011100001001: oled_data = 16'b1000101101101000;
				18'b001010011110001001: oled_data = 16'b1000101110001001;
				18'b001010100000001001: oled_data = 16'b1000101110001010;
				18'b001010100010001001: oled_data = 16'b0101101010101000;
				18'b001010100100001001: oled_data = 16'b0011101000000111;
				18'b001010100110001001: oled_data = 16'b0100001000101000;
				18'b001000011000001010: oled_data = 16'b1011010001101100;
				18'b001000011010001010: oled_data = 16'b1011010001001011;
				18'b001000011100001010: oled_data = 16'b1010110001001011;
				18'b001000011110001010: oled_data = 16'b1010010000101011;
				18'b001000100000001010: oled_data = 16'b1101010111110110;
				18'b001000100010001010: oled_data = 16'b1111011010011011;
				18'b001000100100001010: oled_data = 16'b1101110100110110;
				18'b001000100110001010: oled_data = 16'b1101110011010110;
				18'b001000101000001010: oled_data = 16'b1101110011010101;
				18'b001000101010001010: oled_data = 16'b1101110011010101;
				18'b001000101100001010: oled_data = 16'b1101110011010101;
				18'b001000101110001010: oled_data = 16'b1101110011010101;
				18'b001000110000001010: oled_data = 16'b1101110011010101;
				18'b001000110010001010: oled_data = 16'b1101110011010101;
				18'b001000110100001010: oled_data = 16'b1101110011010110;
				18'b001000110110001010: oled_data = 16'b1101110010010101;
				18'b001000111000001010: oled_data = 16'b1101110010110101;
				18'b001000111010001010: oled_data = 16'b1101110011010101;
				18'b001000111100001010: oled_data = 16'b1101110011010101;
				18'b001000111110001010: oled_data = 16'b1101110011010101;
				18'b001001000000001010: oled_data = 16'b1101110011010101;
				18'b001001000010001010: oled_data = 16'b1101110011010101;
				18'b001001000100001010: oled_data = 16'b1101110011010101;
				18'b001001000110001010: oled_data = 16'b1101110011010101;
				18'b001001001000001010: oled_data = 16'b1101110011010101;
				18'b001001001010001010: oled_data = 16'b1101110011010101;
				18'b001001001100001010: oled_data = 16'b1101110011010101;
				18'b001001001110001010: oled_data = 16'b1101110011010101;
				18'b001001010000001010: oled_data = 16'b1101110011010101;
				18'b001001010010001010: oled_data = 16'b1101110011010101;
				18'b001001010100001010: oled_data = 16'b1101110011010101;
				18'b001001010110001010: oled_data = 16'b1101110011010110;
				18'b001001011000001010: oled_data = 16'b1101010001110100;
				18'b001001011010001010: oled_data = 16'b1101110010110101;
				18'b001001011100001010: oled_data = 16'b1101110011010101;
				18'b001001011110001010: oled_data = 16'b1101110011010101;
				18'b001001100000001010: oled_data = 16'b1101110011010101;
				18'b001001100010001010: oled_data = 16'b1101110011010101;
				18'b001001100100001010: oled_data = 16'b1101110011010101;
				18'b001001100110001010: oled_data = 16'b1101110011010101;
				18'b001001101000001010: oled_data = 16'b1101110011010110;
				18'b001001101010001010: oled_data = 16'b1101010010010100;
				18'b001001101100001010: oled_data = 16'b1101110010110101;
				18'b001001101110001010: oled_data = 16'b1101110011010110;
				18'b001001110000001010: oled_data = 16'b1101110011010110;
				18'b001001110010001010: oled_data = 16'b1101010010010101;
				18'b001001110100001010: oled_data = 16'b1101110010110101;
				18'b001001110110001010: oled_data = 16'b1101110011010110;
				18'b001001111000001010: oled_data = 16'b1101110011010101;
				18'b001001111010001010: oled_data = 16'b1101110011010101;
				18'b001001111100001010: oled_data = 16'b1101010001110100;
				18'b001001111110001010: oled_data = 16'b1101110011010101;
				18'b001010000000001010: oled_data = 16'b1101110011010101;
				18'b001010000010001010: oled_data = 16'b1101110011010101;
				18'b001010000100001010: oled_data = 16'b1101110100010110;
				18'b001010000110001010: oled_data = 16'b1111011010111100;
				18'b001010001000001010: oled_data = 16'b1100010101010101;
				18'b001010001010001010: oled_data = 16'b0011100101100101;
				18'b001010001100001010: oled_data = 16'b0100000111000110;
				18'b001010001110001010: oled_data = 16'b0101001000100110;
				18'b001010010000001010: oled_data = 16'b0101101010000111;
				18'b001010010010001010: oled_data = 16'b0110101011001000;
				18'b001010010100001010: oled_data = 16'b0111101011101000;
				18'b001010010110001010: oled_data = 16'b1000001100101000;
				18'b001010011000001010: oled_data = 16'b1000101101001000;
				18'b001010011010001010: oled_data = 16'b1000101101101000;
				18'b001010011100001010: oled_data = 16'b1000101110001000;
				18'b001010011110001010: oled_data = 16'b1000101110001000;
				18'b001010100000001010: oled_data = 16'b1000101110001001;
				18'b001010100010001010: oled_data = 16'b0111001011101001;
				18'b001010100100001010: oled_data = 16'b1001001101001101;
				18'b001010100110001010: oled_data = 16'b1011010000110001;
				18'b001000011000001011: oled_data = 16'b1001101111001010;
				18'b001000011010001011: oled_data = 16'b1000101110001010;
				18'b001000011100001011: oled_data = 16'b0111001100001001;
				18'b001000011110001011: oled_data = 16'b1000001110101100;
				18'b001000100000001011: oled_data = 16'b1111011010111011;
				18'b001000100010001011: oled_data = 16'b1110010110111000;
				18'b001000100100001011: oled_data = 16'b1101110011010101;
				18'b001000100110001011: oled_data = 16'b1101110011010110;
				18'b001000101000001011: oled_data = 16'b1101110011010101;
				18'b001000101010001011: oled_data = 16'b1101110011010101;
				18'b001000101100001011: oled_data = 16'b1101110011010101;
				18'b001000101110001011: oled_data = 16'b1101110011010101;
				18'b001000110000001011: oled_data = 16'b1101110011010101;
				18'b001000110010001011: oled_data = 16'b1101110011010101;
				18'b001000110100001011: oled_data = 16'b1101110010110101;
				18'b001000110110001011: oled_data = 16'b1101010001110100;
				18'b001000111000001011: oled_data = 16'b1101110011010101;
				18'b001000111010001011: oled_data = 16'b1101110011010101;
				18'b001000111100001011: oled_data = 16'b1101110011010101;
				18'b001000111110001011: oled_data = 16'b1101110011010101;
				18'b001001000000001011: oled_data = 16'b1101110011010101;
				18'b001001000010001011: oled_data = 16'b1101110011010101;
				18'b001001000100001011: oled_data = 16'b1101110011010101;
				18'b001001000110001011: oled_data = 16'b1101110011010101;
				18'b001001001000001011: oled_data = 16'b1101110011010101;
				18'b001001001010001011: oled_data = 16'b1101110011010101;
				18'b001001001100001011: oled_data = 16'b1101110011010101;
				18'b001001001110001011: oled_data = 16'b1101110011010101;
				18'b001001010000001011: oled_data = 16'b1101110011010101;
				18'b001001010010001011: oled_data = 16'b1101110011010101;
				18'b001001010100001011: oled_data = 16'b1101110011010110;
				18'b001001010110001011: oled_data = 16'b1101110011010110;
				18'b001001011000001011: oled_data = 16'b1101010001110100;
				18'b001001011010001011: oled_data = 16'b1101110011010101;
				18'b001001011100001011: oled_data = 16'b1101110011010101;
				18'b001001011110001011: oled_data = 16'b1101110011010101;
				18'b001001100000001011: oled_data = 16'b1101110011010101;
				18'b001001100010001011: oled_data = 16'b1101110011010101;
				18'b001001100100001011: oled_data = 16'b1101110011010101;
				18'b001001100110001011: oled_data = 16'b1101110011010101;
				18'b001001101000001011: oled_data = 16'b1101110011010101;
				18'b001001101010001011: oled_data = 16'b1101110010110101;
				18'b001001101100001011: oled_data = 16'b1101010010010100;
				18'b001001101110001011: oled_data = 16'b1101110011010110;
				18'b001001110000001011: oled_data = 16'b1101110011010101;
				18'b001001110010001011: oled_data = 16'b1101110010110101;
				18'b001001110100001011: oled_data = 16'b1101010001110100;
				18'b001001110110001011: oled_data = 16'b1101110011010110;
				18'b001001111000001011: oled_data = 16'b1101110011010101;
				18'b001001111010001011: oled_data = 16'b1110010010110101;
				18'b001001111100001011: oled_data = 16'b1101110010010101;
				18'b001001111110001011: oled_data = 16'b1101110010110101;
				18'b001010000000001011: oled_data = 16'b1101110011010101;
				18'b001010000010001011: oled_data = 16'b1101110011010101;
				18'b001010000100001011: oled_data = 16'b1101010011010101;
				18'b001010000110001011: oled_data = 16'b1110011000111001;
				18'b001010001000001011: oled_data = 16'b1110111010111011;
				18'b001010001010001011: oled_data = 16'b0100000111101000;
				18'b001010001100001011: oled_data = 16'b0001100100000101;
				18'b001010001110001011: oled_data = 16'b0010000101000101;
				18'b001010010000001011: oled_data = 16'b0010000101100110;
				18'b001010010010001011: oled_data = 16'b0010100110000111;
				18'b001010010100001011: oled_data = 16'b0011100111000111;
				18'b001010010110001011: oled_data = 16'b0100001000000111;
				18'b001010011000001011: oled_data = 16'b0101001000100111;
				18'b001010011010001011: oled_data = 16'b0101101001100111;
				18'b001010011100001011: oled_data = 16'b0111001011001000;
				18'b001010011110001011: oled_data = 16'b1010001110001100;
				18'b001010100000001011: oled_data = 16'b1100010001010000;
				18'b001010100010001011: oled_data = 16'b1101110010110010;
				18'b001010100100001011: oled_data = 16'b1101110001010001;
				18'b001010100110001011: oled_data = 16'b1100101110001110;
				18'b001000011000001100: oled_data = 16'b0101101010101000;
				18'b001000011010001100: oled_data = 16'b0110001010101001;
				18'b001000011100001100: oled_data = 16'b0110101010101001;
				18'b001000011110001100: oled_data = 16'b1010110011010001;
				18'b001000100000001100: oled_data = 16'b1111111010111100;
				18'b001000100010001100: oled_data = 16'b1110010100010110;
				18'b001000100100001100: oled_data = 16'b1110010011010101;
				18'b001000100110001100: oled_data = 16'b1101110011010101;
				18'b001000101000001100: oled_data = 16'b1101110011010101;
				18'b001000101010001100: oled_data = 16'b1101110011010101;
				18'b001000101100001100: oled_data = 16'b1101110011010101;
				18'b001000101110001100: oled_data = 16'b1101110011010101;
				18'b001000110000001100: oled_data = 16'b1101110011010101;
				18'b001000110010001100: oled_data = 16'b1101110011010101;
				18'b001000110100001100: oled_data = 16'b1101010001110100;
				18'b001000110110001100: oled_data = 16'b1101110011010110;
				18'b001000111000001100: oled_data = 16'b1101110011010110;
				18'b001000111010001100: oled_data = 16'b1101110011010101;
				18'b001000111100001100: oled_data = 16'b1101110011010101;
				18'b001000111110001100: oled_data = 16'b1101110011010101;
				18'b001001000000001100: oled_data = 16'b1101110011010101;
				18'b001001000010001100: oled_data = 16'b1101110011010101;
				18'b001001000100001100: oled_data = 16'b1101110011010101;
				18'b001001000110001100: oled_data = 16'b1101110011010101;
				18'b001001001000001100: oled_data = 16'b1101110011010101;
				18'b001001001010001100: oled_data = 16'b1101110011010101;
				18'b001001001100001100: oled_data = 16'b1101110011010101;
				18'b001001001110001100: oled_data = 16'b1101110011010101;
				18'b001001010000001100: oled_data = 16'b1101110011010101;
				18'b001001010010001100: oled_data = 16'b1101110011010101;
				18'b001001010100001100: oled_data = 16'b1101110011010101;
				18'b001001010110001100: oled_data = 16'b1101110010110101;
				18'b001001011000001100: oled_data = 16'b1101010001110100;
				18'b001001011010001100: oled_data = 16'b1101110011010110;
				18'b001001011100001100: oled_data = 16'b1101110011010101;
				18'b001001011110001100: oled_data = 16'b1101110011010101;
				18'b001001100000001100: oled_data = 16'b1101110011110110;
				18'b001001100010001100: oled_data = 16'b1101110011010101;
				18'b001001100100001100: oled_data = 16'b1101110011010101;
				18'b001001100110001100: oled_data = 16'b1101110011010101;
				18'b001001101000001100: oled_data = 16'b1101110011010101;
				18'b001001101010001100: oled_data = 16'b1101110011010101;
				18'b001001101100001100: oled_data = 16'b1101010010010100;
				18'b001001101110001100: oled_data = 16'b1101110011010110;
				18'b001001110000001100: oled_data = 16'b1101110011010101;
				18'b001001110010001100: oled_data = 16'b1101110011010101;
				18'b001001110100001100: oled_data = 16'b1101010001110100;
				18'b001001110110001100: oled_data = 16'b1101110011010101;
				18'b001001111000001100: oled_data = 16'b1101110011010101;
				18'b001001111010001100: oled_data = 16'b1110010011010110;
				18'b001001111100001100: oled_data = 16'b1101110010010101;
				18'b001001111110001100: oled_data = 16'b1101010010010101;
				18'b001010000000001100: oled_data = 16'b1101110011010110;
				18'b001010000010001100: oled_data = 16'b1101110011010101;
				18'b001010000100001100: oled_data = 16'b1101110011010101;
				18'b001010000110001100: oled_data = 16'b1101110101010111;
				18'b001010001000001100: oled_data = 16'b1111111011111100;
				18'b001010001010001100: oled_data = 16'b0111001100101101;
				18'b001010001100001100: oled_data = 16'b0001100011100100;
				18'b001010001110001100: oled_data = 16'b0010000101000101;
				18'b001010010000001100: oled_data = 16'b0010000101000110;
				18'b001010010010001100: oled_data = 16'b0010100101100110;
				18'b001010010100001100: oled_data = 16'b0010100110000111;
				18'b001010010110001100: oled_data = 16'b0010100110000111;
				18'b001010011000001100: oled_data = 16'b0010100110100111;
				18'b001010011010001100: oled_data = 16'b0110101010101010;
				18'b001010011100001100: oled_data = 16'b1011110001010001;
				18'b001010011110001100: oled_data = 16'b1110010011010100;
				18'b001010100000001100: oled_data = 16'b1101110000110001;
				18'b001010100010001100: oled_data = 16'b1100001100001100;
				18'b001010100100001100: oled_data = 16'b1010101001001001;
				18'b001010100110001100: oled_data = 16'b1010101000001000;
				18'b001000011000001101: oled_data = 16'b1001110000001011;
				18'b001000011010001101: oled_data = 16'b1001010010110000;
				18'b001000011100001101: oled_data = 16'b1000110100110011;
				18'b001000011110001101: oled_data = 16'b1001111000010111;
				18'b001000100000001101: oled_data = 16'b1011011000011001;
				18'b001000100010001101: oled_data = 16'b1100010100010111;
				18'b001000100100001101: oled_data = 16'b1101110011010110;
				18'b001000100110001101: oled_data = 16'b1110010011010101;
				18'b001000101000001101: oled_data = 16'b1101110011010101;
				18'b001000101010001101: oled_data = 16'b1101110011010101;
				18'b001000101100001101: oled_data = 16'b1101110011010101;
				18'b001000101110001101: oled_data = 16'b1101110011010101;
				18'b001000110000001101: oled_data = 16'b1101110011010110;
				18'b001000110010001101: oled_data = 16'b1101010001110100;
				18'b001000110100001101: oled_data = 16'b1101110010110101;
				18'b001000110110001101: oled_data = 16'b1110010011110110;
				18'b001000111000001101: oled_data = 16'b1101110011010101;
				18'b001000111010001101: oled_data = 16'b1110010011110110;
				18'b001000111100001101: oled_data = 16'b1110010011110110;
				18'b001000111110001101: oled_data = 16'b1101110011010101;
				18'b001001000000001101: oled_data = 16'b1101110011010101;
				18'b001001000010001101: oled_data = 16'b1101110011010101;
				18'b001001000100001101: oled_data = 16'b1101110011010101;
				18'b001001000110001101: oled_data = 16'b1101110011010101;
				18'b001001001000001101: oled_data = 16'b1101110011010101;
				18'b001001001010001101: oled_data = 16'b1101110011010101;
				18'b001001001100001101: oled_data = 16'b1101110011010101;
				18'b001001001110001101: oled_data = 16'b1101110011010101;
				18'b001001010000001101: oled_data = 16'b1101110011010101;
				18'b001001010010001101: oled_data = 16'b1101110011010101;
				18'b001001010100001101: oled_data = 16'b1101110011010101;
				18'b001001010110001101: oled_data = 16'b1101110010110101;
				18'b001001011000001101: oled_data = 16'b1101010010010100;
				18'b001001011010001101: oled_data = 16'b1101110011010110;
				18'b001001011100001101: oled_data = 16'b1101110011010101;
				18'b001001011110001101: oled_data = 16'b1101110011010110;
				18'b001001100000001101: oled_data = 16'b1110110101111000;
				18'b001001100010001101: oled_data = 16'b1101110011010101;
				18'b001001100100001101: oled_data = 16'b1101110011010101;
				18'b001001100110001101: oled_data = 16'b1101110011010101;
				18'b001001101000001101: oled_data = 16'b1101110011010101;
				18'b001001101010001101: oled_data = 16'b1101110011010101;
				18'b001001101100001101: oled_data = 16'b1101010001110100;
				18'b001001101110001101: oled_data = 16'b1101110011010101;
				18'b001001110000001101: oled_data = 16'b1101110011010101;
				18'b001001110010001101: oled_data = 16'b1101110011010110;
				18'b001001110100001101: oled_data = 16'b1101010001110100;
				18'b001001110110001101: oled_data = 16'b1101110010110101;
				18'b001001111000001101: oled_data = 16'b1101110011010101;
				18'b001001111010001101: oled_data = 16'b1101110011010101;
				18'b001001111100001101: oled_data = 16'b1101110010110101;
				18'b001001111110001101: oled_data = 16'b1101010010010100;
				18'b001010000000001101: oled_data = 16'b1101110011010110;
				18'b001010000010001101: oled_data = 16'b1101110011010101;
				18'b001010000100001101: oled_data = 16'b1101110011010101;
				18'b001010000110001101: oled_data = 16'b1101010011110110;
				18'b001010001000001101: oled_data = 16'b1111011011011011;
				18'b001010001010001101: oled_data = 16'b1010010010110011;
				18'b001010001100001101: oled_data = 16'b0001100011100100;
				18'b001010001110001101: oled_data = 16'b0010000100100101;
				18'b001010010000001101: oled_data = 16'b0010000101000110;
				18'b001010010010001101: oled_data = 16'b0010000101100110;
				18'b001010010100001101: oled_data = 16'b0010000101000110;
				18'b001010010110001101: oled_data = 16'b0100001000001000;
				18'b001010011000001101: oled_data = 16'b1010101111110000;
				18'b001010011010001101: oled_data = 16'b1110010100010100;
				18'b001010011100001101: oled_data = 16'b1110010010010010;
				18'b001010011110001101: oled_data = 16'b1100001100101101;
				18'b001010100000001101: oled_data = 16'b1011001001001001;
				18'b001010100010001101: oled_data = 16'b1011001000101000;
				18'b001010100100001101: oled_data = 16'b1010101000101000;
				18'b001010100110001101: oled_data = 16'b1010101000001000;
				18'b001000011000001110: oled_data = 16'b1001010011001111;
				18'b001000011010001110: oled_data = 16'b1000111000111001;
				18'b001000011100001110: oled_data = 16'b1010111100011101;
				18'b001000011110001110: oled_data = 16'b1010111011111100;
				18'b001000100000001110: oled_data = 16'b1000111010011010;
				18'b001000100010001110: oled_data = 16'b1000011000111010;
				18'b001000100100001110: oled_data = 16'b1000110111011001;
				18'b001000100110001110: oled_data = 16'b1011010100010110;
				18'b001000101000001110: oled_data = 16'b1101110010110101;
				18'b001000101010001110: oled_data = 16'b1101110011010101;
				18'b001000101100001110: oled_data = 16'b1101110011010101;
				18'b001000101110001110: oled_data = 16'b1101110011010101;
				18'b001000110000001110: oled_data = 16'b1101110010110101;
				18'b001000110010001110: oled_data = 16'b1101010001110100;
				18'b001000110100001110: oled_data = 16'b1101110011010101;
				18'b001000110110001110: oled_data = 16'b1101110011010101;
				18'b001000111000001110: oled_data = 16'b1101110011010110;
				18'b001000111010001110: oled_data = 16'b1110110100110111;
				18'b001000111100001110: oled_data = 16'b1110010011010110;
				18'b001000111110001110: oled_data = 16'b1101110011010101;
				18'b001001000000001110: oled_data = 16'b1101110011010101;
				18'b001001000010001110: oled_data = 16'b1101110011010101;
				18'b001001000100001110: oled_data = 16'b1101110011010110;
				18'b001001000110001110: oled_data = 16'b1101110010010101;
				18'b001001001000001110: oled_data = 16'b1101010001110100;
				18'b001001001010001110: oled_data = 16'b1101110011010110;
				18'b001001001100001110: oled_data = 16'b1101110011010101;
				18'b001001001110001110: oled_data = 16'b1101110011010101;
				18'b001001010000001110: oled_data = 16'b1101110011010101;
				18'b001001010010001110: oled_data = 16'b1101110011010101;
				18'b001001010100001110: oled_data = 16'b1101110011010110;
				18'b001001010110001110: oled_data = 16'b1101110010010101;
				18'b001001011000001110: oled_data = 16'b1101110010010101;
				18'b001001011010001110: oled_data = 16'b1101110011010110;
				18'b001001011100001110: oled_data = 16'b1101110011010101;
				18'b001001011110001110: oled_data = 16'b1110010011110110;
				18'b001001100000001110: oled_data = 16'b1110110110011000;
				18'b001001100010001110: oled_data = 16'b1101110011010101;
				18'b001001100100001110: oled_data = 16'b1101110011010101;
				18'b001001100110001110: oled_data = 16'b1101110011010101;
				18'b001001101000001110: oled_data = 16'b1101110011010101;
				18'b001001101010001110: oled_data = 16'b1101110011010110;
				18'b001001101100001110: oled_data = 16'b1101010001110100;
				18'b001001101110001110: oled_data = 16'b1101110011010101;
				18'b001001110000001110: oled_data = 16'b1101110011010101;
				18'b001001110010001110: oled_data = 16'b1101110011010110;
				18'b001001110100001110: oled_data = 16'b1101010010010100;
				18'b001001110110001110: oled_data = 16'b1101110010110101;
				18'b001001111000001110: oled_data = 16'b1101110011010101;
				18'b001001111010001110: oled_data = 16'b1101110011010101;
				18'b001001111100001110: oled_data = 16'b1101110011010101;
				18'b001001111110001110: oled_data = 16'b1101010001110100;
				18'b001010000000001110: oled_data = 16'b1101110011010101;
				18'b001010000010001110: oled_data = 16'b1101110011010101;
				18'b001010000100001110: oled_data = 16'b1101110010010101;
				18'b001010000110001110: oled_data = 16'b1101110011010101;
				18'b001010001000001110: oled_data = 16'b1110111000111010;
				18'b001010001010001110: oled_data = 16'b1100110110110111;
				18'b001010001100001110: oled_data = 16'b0010000100100101;
				18'b001010001110001110: oled_data = 16'b0001100100100101;
				18'b001010010000001110: oled_data = 16'b0010000101000110;
				18'b001010010010001110: oled_data = 16'b0010000101000101;
				18'b001010010100001110: oled_data = 16'b0110001010001010;
				18'b001010010110001110: oled_data = 16'b1101010010010010;
				18'b001010011000001110: oled_data = 16'b1110110011110100;
				18'b001010011010001110: oled_data = 16'b1101001111001111;
				18'b001010011100001110: oled_data = 16'b1011101010001010;
				18'b001010011110001110: oled_data = 16'b1011001000001000;
				18'b001010100000001110: oled_data = 16'b1011001000101001;
				18'b001010100010001110: oled_data = 16'b1011001000101000;
				18'b001010100100001110: oled_data = 16'b1010101000101000;
				18'b001010100110001110: oled_data = 16'b1010101000001000;
				18'b001000011000001111: oled_data = 16'b1000010101110101;
				18'b001000011010001111: oled_data = 16'b1001011010011011;
				18'b001000011100001111: oled_data = 16'b1011011100111100;
				18'b001000011110001111: oled_data = 16'b1011111100111101;
				18'b001000100000001111: oled_data = 16'b1011011100011100;
				18'b001000100010001111: oled_data = 16'b0111010110111001;
				18'b001000100100001111: oled_data = 16'b0111011000011010;
				18'b001000100110001111: oled_data = 16'b0111111000011010;
				18'b001000101000001111: oled_data = 16'b1011110100010110;
				18'b001000101010001111: oled_data = 16'b1110010011010101;
				18'b001000101100001111: oled_data = 16'b1101110011010101;
				18'b001000101110001111: oled_data = 16'b1101110011010110;
				18'b001000110000001111: oled_data = 16'b1101010010010100;
				18'b001000110010001111: oled_data = 16'b1101110011010101;
				18'b001000110100001111: oled_data = 16'b1101110011010101;
				18'b001000110110001111: oled_data = 16'b1101110011010101;
				18'b001000111000001111: oled_data = 16'b1110010011110110;
				18'b001000111010001111: oled_data = 16'b1110010011110110;
				18'b001000111100001111: oled_data = 16'b1101110011010101;
				18'b001000111110001111: oled_data = 16'b1101110011010101;
				18'b001001000000001111: oled_data = 16'b1101110011010101;
				18'b001001000010001111: oled_data = 16'b1101110011010101;
				18'b001001000100001111: oled_data = 16'b1101110011010110;
				18'b001001000110001111: oled_data = 16'b1101010001010100;
				18'b001001001000001111: oled_data = 16'b1101110010110101;
				18'b001001001010001111: oled_data = 16'b1101110011010110;
				18'b001001001100001111: oled_data = 16'b1101110011010101;
				18'b001001001110001111: oled_data = 16'b1101110010110101;
				18'b001001010000001111: oled_data = 16'b1101110010110101;
				18'b001001010010001111: oled_data = 16'b1101110011010110;
				18'b001001010100001111: oled_data = 16'b1101110011010110;
				18'b001001010110001111: oled_data = 16'b1101010010010100;
				18'b001001011000001111: oled_data = 16'b1101110010110101;
				18'b001001011010001111: oled_data = 16'b1101110011010101;
				18'b001001011100001111: oled_data = 16'b1101110011010101;
				18'b001001011110001111: oled_data = 16'b1110010011110110;
				18'b001001100000001111: oled_data = 16'b1110010101010111;
				18'b001001100010001111: oled_data = 16'b1101110010110101;
				18'b001001100100001111: oled_data = 16'b1101110011010101;
				18'b001001100110001111: oled_data = 16'b1101110011010101;
				18'b001001101000001111: oled_data = 16'b1101110011010101;
				18'b001001101010001111: oled_data = 16'b1101110011010110;
				18'b001001101100001111: oled_data = 16'b1101010010010100;
				18'b001001101110001111: oled_data = 16'b1101110010110101;
				18'b001001110000001111: oled_data = 16'b1101110011010101;
				18'b001001110010001111: oled_data = 16'b1101110011010110;
				18'b001001110100001111: oled_data = 16'b1101010010010100;
				18'b001001110110001111: oled_data = 16'b1101110010010101;
				18'b001001111000001111: oled_data = 16'b1101110011010110;
				18'b001001111010001111: oled_data = 16'b1101110011010101;
				18'b001001111100001111: oled_data = 16'b1101110011010101;
				18'b001001111110001111: oled_data = 16'b1101010001110100;
				18'b001010000000001111: oled_data = 16'b1101110011010101;
				18'b001010000010001111: oled_data = 16'b1101110011010110;
				18'b001010000100001111: oled_data = 16'b1101010010010100;
				18'b001010000110001111: oled_data = 16'b1101110010110101;
				18'b001010001000001111: oled_data = 16'b1101110110111000;
				18'b001010001010001111: oled_data = 16'b1110011001111010;
				18'b001010001100001111: oled_data = 16'b0011000110100111;
				18'b001010001110001111: oled_data = 16'b0001000100100100;
				18'b001010010000001111: oled_data = 16'b0001100100100101;
				18'b001010010010001111: oled_data = 16'b0111101100001100;
				18'b001010010100001111: oled_data = 16'b1110010100010100;
				18'b001010010110001111: oled_data = 16'b1110010010110010;
				18'b001010011000001111: oled_data = 16'b1100001100001100;
				18'b001010011010001111: oled_data = 16'b1011001000101001;
				18'b001010011100001111: oled_data = 16'b1011001000101001;
				18'b001010011110001111: oled_data = 16'b1011001000101001;
				18'b001010100000001111: oled_data = 16'b1011001000101001;
				18'b001010100010001111: oled_data = 16'b1011001000101000;
				18'b001010100100001111: oled_data = 16'b1010101000101000;
				18'b001010100110001111: oled_data = 16'b1010101000001000;
				18'b001000011000010000: oled_data = 16'b0111011000011010;
				18'b001000011010010000: oled_data = 16'b1001011010011011;
				18'b001000011100010000: oled_data = 16'b1011011101011100;
				18'b001000011110010000: oled_data = 16'b1001111001111011;
				18'b001000100000010000: oled_data = 16'b0111010100110111;
				18'b001000100010010000: oled_data = 16'b0100110001110110;
				18'b001000100100010000: oled_data = 16'b0101010010010110;
				18'b001000100110010000: oled_data = 16'b0111011000011010;
				18'b001000101000010000: oled_data = 16'b1010010101111000;
				18'b001000101010010000: oled_data = 16'b1110010010110101;
				18'b001000101100010000: oled_data = 16'b1101110011010110;
				18'b001000101110010000: oled_data = 16'b1101010010010101;
				18'b001000110000010000: oled_data = 16'b1101110010010101;
				18'b001000110010010000: oled_data = 16'b1110010011010110;
				18'b001000110100010000: oled_data = 16'b1101110011010101;
				18'b001000110110010000: oled_data = 16'b1101110011010101;
				18'b001000111000010000: oled_data = 16'b1101110011010110;
				18'b001000111010010000: oled_data = 16'b1101110011010110;
				18'b001000111100010000: oled_data = 16'b1101110011010101;
				18'b001000111110010000: oled_data = 16'b1101110011010101;
				18'b001001000000010000: oled_data = 16'b1101110011010101;
				18'b001001000010010000: oled_data = 16'b1101110011010101;
				18'b001001000100010000: oled_data = 16'b1101110010110101;
				18'b001001000110010000: oled_data = 16'b1101010001110100;
				18'b001001001000010000: oled_data = 16'b1101110011010110;
				18'b001001001010010000: oled_data = 16'b1101110011010110;
				18'b001001001100010000: oled_data = 16'b1101110011010110;
				18'b001001001110010000: oled_data = 16'b1101010010010100;
				18'b001001010000010000: oled_data = 16'b1101110010110101;
				18'b001001010010010000: oled_data = 16'b1101110011010101;
				18'b001001010100010000: oled_data = 16'b1101110011010110;
				18'b001001010110010000: oled_data = 16'b1101010001110100;
				18'b001001011000010000: oled_data = 16'b1101110010110101;
				18'b001001011010010000: oled_data = 16'b1101110011010101;
				18'b001001011100010000: oled_data = 16'b1101110011010101;
				18'b001001011110010000: oled_data = 16'b1101110011110110;
				18'b001001100000010000: oled_data = 16'b1110010100010110;
				18'b001001100010010000: oled_data = 16'b1101110011010101;
				18'b001001100100010000: oled_data = 16'b1101110011010101;
				18'b001001100110010000: oled_data = 16'b1101110011010101;
				18'b001001101000010000: oled_data = 16'b1101110011010101;
				18'b001001101010010000: oled_data = 16'b1101110011010110;
				18'b001001101100010000: oled_data = 16'b1101010010010100;
				18'b001001101110010000: oled_data = 16'b1101110010110101;
				18'b001001110000010000: oled_data = 16'b1101110011010101;
				18'b001001110010010000: oled_data = 16'b1101110011010110;
				18'b001001110100010000: oled_data = 16'b1101010010010100;
				18'b001001110110010000: oled_data = 16'b1101010001110100;
				18'b001001111000010000: oled_data = 16'b1101110011010110;
				18'b001001111010010000: oled_data = 16'b1101110011010101;
				18'b001001111100010000: oled_data = 16'b1101110011010101;
				18'b001001111110010000: oled_data = 16'b1101010001110100;
				18'b001010000000010000: oled_data = 16'b1101110011010101;
				18'b001010000010010000: oled_data = 16'b1101110011010101;
				18'b001010000100010000: oled_data = 16'b1101110010110101;
				18'b001010000110010000: oled_data = 16'b1101010010010101;
				18'b001010001000010000: oled_data = 16'b1101110101110111;
				18'b001010001010010000: oled_data = 16'b1110111011011011;
				18'b001010001100010000: oled_data = 16'b0100001000101001;
				18'b001010001110010000: oled_data = 16'b0001100011100100;
				18'b001010010000010000: oled_data = 16'b1000101100101110;
				18'b001010010010010000: oled_data = 16'b1110110100010101;
				18'b001010010100010000: oled_data = 16'b1101110001010001;
				18'b001010010110010000: oled_data = 16'b1011101010101010;
				18'b001010011000010000: oled_data = 16'b1011001000101001;
				18'b001010011010010000: oled_data = 16'b1011001000101001;
				18'b001010011100010000: oled_data = 16'b1011001000101001;
				18'b001010011110010000: oled_data = 16'b1011001000101001;
				18'b001010100000010000: oled_data = 16'b1011001000101001;
				18'b001010100010010000: oled_data = 16'b1011001000101000;
				18'b001010100100010000: oled_data = 16'b1010101000101000;
				18'b001010100110010000: oled_data = 16'b1010101000001000;
				18'b001000011000010001: oled_data = 16'b0111011000011010;
				18'b001000011010010001: oled_data = 16'b1000011000111010;
				18'b001000011100010001: oled_data = 16'b1001011010011011;
				18'b001000011110010001: oled_data = 16'b0101010010010110;
				18'b001000100000010001: oled_data = 16'b0100010001010110;
				18'b001000100010010001: oled_data = 16'b0100110001010110;
				18'b001000100100010001: oled_data = 16'b0100110001010101;
				18'b001000100110010001: oled_data = 16'b0110010110011001;
				18'b001000101000010001: oled_data = 16'b1010010101111000;
				18'b001000101010010001: oled_data = 16'b1110010010110110;
				18'b001000101100010001: oled_data = 16'b1101110011010101;
				18'b001000101110010001: oled_data = 16'b1101010001110100;
				18'b001000110000010001: oled_data = 16'b1101110011010110;
				18'b001000110010010001: oled_data = 16'b1101110011010101;
				18'b001000110100010001: oled_data = 16'b1101110011010101;
				18'b001000110110010001: oled_data = 16'b1101110010110101;
				18'b001000111000010001: oled_data = 16'b1101110011010101;
				18'b001000111010010001: oled_data = 16'b1101110011010101;
				18'b001000111100010001: oled_data = 16'b1101110011010101;
				18'b001000111110010001: oled_data = 16'b1101110011010101;
				18'b001001000000010001: oled_data = 16'b1101110011010101;
				18'b001001000010010001: oled_data = 16'b1101110011010110;
				18'b001001000100010001: oled_data = 16'b1101010001110100;
				18'b001001000110010001: oled_data = 16'b1101110010110101;
				18'b001001001000010001: oled_data = 16'b1101110011010101;
				18'b001001001010010001: oled_data = 16'b1101110011010101;
				18'b001001001100010001: oled_data = 16'b1101110011010110;
				18'b001001001110010001: oled_data = 16'b1101010001110100;
				18'b001001010000010001: oled_data = 16'b1101110010110101;
				18'b001001010010010001: oled_data = 16'b1101110011010101;
				18'b001001010100010001: oled_data = 16'b1101110011010110;
				18'b001001010110010001: oled_data = 16'b1101010001110100;
				18'b001001011000010001: oled_data = 16'b1101110010110101;
				18'b001001011010010001: oled_data = 16'b1101110011010101;
				18'b001001011100010001: oled_data = 16'b1101110011010101;
				18'b001001011110010001: oled_data = 16'b1101110011010101;
				18'b001001100000010001: oled_data = 16'b1101110011010101;
				18'b001001100010010001: oled_data = 16'b1101110011010101;
				18'b001001100100010001: oled_data = 16'b1101110011010101;
				18'b001001100110010001: oled_data = 16'b1101110011010101;
				18'b001001101000010001: oled_data = 16'b1101110011010101;
				18'b001001101010010001: oled_data = 16'b1101110011010110;
				18'b001001101100010001: oled_data = 16'b1101010001110100;
				18'b001001101110010001: oled_data = 16'b1101110010110101;
				18'b001001110000010001: oled_data = 16'b1101110011010110;
				18'b001001110010010001: oled_data = 16'b1101110011010110;
				18'b001001110100010001: oled_data = 16'b1101010010010100;
				18'b001001110110010001: oled_data = 16'b1101010001110100;
				18'b001001111000010001: oled_data = 16'b1101110011010110;
				18'b001001111010010001: oled_data = 16'b1101110011010101;
				18'b001001111100010001: oled_data = 16'b1101110011010101;
				18'b001001111110010001: oled_data = 16'b1100110000110011;
				18'b001010000000010001: oled_data = 16'b1101110011010101;
				18'b001010000010010001: oled_data = 16'b1101110011010101;
				18'b001010000100010001: oled_data = 16'b1101110010110101;
				18'b001010000110010001: oled_data = 16'b1101010010010100;
				18'b001010001000010001: oled_data = 16'b1101010100010110;
				18'b001010001010010001: oled_data = 16'b1110111010111011;
				18'b001010001100010001: oled_data = 16'b0101001010001011;
				18'b001010001110010001: oled_data = 16'b1000001011101100;
				18'b001010010000010001: oled_data = 16'b1110110100110101;
				18'b001010010010010001: oled_data = 16'b1101110000010000;
				18'b001010010100010001: oled_data = 16'b1011001010001010;
				18'b001010010110010001: oled_data = 16'b1011001000101001;
				18'b001010011000010001: oled_data = 16'b1011001001001001;
				18'b001010011010010001: oled_data = 16'b1011001000101001;
				18'b001010011100010001: oled_data = 16'b1011001001001001;
				18'b001010011110010001: oled_data = 16'b1011001000101001;
				18'b001010100000010001: oled_data = 16'b1011001000101001;
				18'b001010100010010001: oled_data = 16'b1011001000101000;
				18'b001010100100010001: oled_data = 16'b1011001000001000;
				18'b001010100110010001: oled_data = 16'b1011001000001000;
				18'b001000011000010010: oled_data = 16'b0111011000011010;
				18'b001000011010010010: oled_data = 16'b0110110110011000;
				18'b001000011100010010: oled_data = 16'b0110110101011000;
				18'b001000011110010010: oled_data = 16'b0100010001010110;
				18'b001000100000010010: oled_data = 16'b0100110001110110;
				18'b001000100010010010: oled_data = 16'b0100110001010110;
				18'b001000100100010010: oled_data = 16'b0100110001010101;
				18'b001000100110010010: oled_data = 16'b0101110101011000;
				18'b001000101000010010: oled_data = 16'b1010010101010111;
				18'b001000101010010010: oled_data = 16'b1110010011010110;
				18'b001000101100010010: oled_data = 16'b1101010010010100;
				18'b001000101110010010: oled_data = 16'b1101110010010101;
				18'b001000110000010010: oled_data = 16'b1101110011010110;
				18'b001000110010010010: oled_data = 16'b1101110011010110;
				18'b001000110100010010: oled_data = 16'b1101110010010101;
				18'b001000110110010010: oled_data = 16'b1101010010010101;
				18'b001000111000010010: oled_data = 16'b1101110011010110;
				18'b001000111010010010: oled_data = 16'b1101110011010101;
				18'b001000111100010010: oled_data = 16'b1101110011010101;
				18'b001000111110010010: oled_data = 16'b1101110011010101;
				18'b001001000000010010: oled_data = 16'b1101110011010101;
				18'b001001000010010010: oled_data = 16'b1101110011010101;
				18'b001001000100010010: oled_data = 16'b1101010010010100;
				18'b001001000110010010: oled_data = 16'b1101110011010101;
				18'b001001001000010010: oled_data = 16'b1101110011010101;
				18'b001001001010010010: oled_data = 16'b1101110011010101;
				18'b001001001100010010: oled_data = 16'b1101110011010101;
				18'b001001001110010010: oled_data = 16'b1101010001110100;
				18'b001001010000010010: oled_data = 16'b1101110011010101;
				18'b001001010010010010: oled_data = 16'b1101110011010101;
				18'b001001010100010010: oled_data = 16'b1101110011010110;
				18'b001001010110010010: oled_data = 16'b1101010010010100;
				18'b001001011000010010: oled_data = 16'b1101110011010101;
				18'b001001011010010010: oled_data = 16'b1101110011010101;
				18'b001001011100010010: oled_data = 16'b1101110011010101;
				18'b001001011110010010: oled_data = 16'b1101110011010101;
				18'b001001100000010010: oled_data = 16'b1101110011010101;
				18'b001001100010010010: oled_data = 16'b1101110011010101;
				18'b001001100100010010: oled_data = 16'b1101110011010101;
				18'b001001100110010010: oled_data = 16'b1101110011010101;
				18'b001001101000010010: oled_data = 16'b1101110011010101;
				18'b001001101010010010: oled_data = 16'b1101110011010110;
				18'b001001101100010010: oled_data = 16'b1101010001110100;
				18'b001001101110010010: oled_data = 16'b1101110010110101;
				18'b001001110000010010: oled_data = 16'b1110010011010110;
				18'b001001110010010010: oled_data = 16'b1101110011010110;
				18'b001001110100010010: oled_data = 16'b1101010010010101;
				18'b001001110110010010: oled_data = 16'b1101010001110100;
				18'b001001111000010010: oled_data = 16'b1101110011010110;
				18'b001001111010010010: oled_data = 16'b1101110011010101;
				18'b001001111100010010: oled_data = 16'b1101110011010110;
				18'b001001111110010010: oled_data = 16'b1100001111110010;
				18'b001010000000010010: oled_data = 16'b1101110010110101;
				18'b001010000010010010: oled_data = 16'b1101110011010101;
				18'b001010000100010010: oled_data = 16'b1101110011010101;
				18'b001010000110010010: oled_data = 16'b1101010001110100;
				18'b001010001000010010: oled_data = 16'b1101010011110101;
				18'b001010001010010010: oled_data = 16'b1110111001011010;
				18'b001010001100010010: oled_data = 16'b1011010001010010;
				18'b001010001110010010: oled_data = 16'b1110010011110100;
				18'b001010010000010010: oled_data = 16'b1101110000110000;
				18'b001010010010010010: oled_data = 16'b1011001001101010;
				18'b001010010100010010: oled_data = 16'b1011001001001001;
				18'b001010010110010010: oled_data = 16'b1011001001001001;
				18'b001010011000010010: oled_data = 16'b1011001001001001;
				18'b001010011010010010: oled_data = 16'b1011001000101001;
				18'b001010011100010010: oled_data = 16'b1011001001001001;
				18'b001010011110010010: oled_data = 16'b1011001000101001;
				18'b001010100000010010: oled_data = 16'b1011001000101001;
				18'b001010100010010010: oled_data = 16'b1011001000101000;
				18'b001010100100010010: oled_data = 16'b1011001000101000;
				18'b001010100110010010: oled_data = 16'b1011001000001000;
				18'b001000011000010011: oled_data = 16'b0111010111111010;
				18'b001000011010010011: oled_data = 16'b0101110100010111;
				18'b001000011100010011: oled_data = 16'b0101110011010111;
				18'b001000011110010011: oled_data = 16'b0100110001010110;
				18'b001000100000010011: oled_data = 16'b0100110001010110;
				18'b001000100010010011: oled_data = 16'b0100110001010101;
				18'b001000100100010011: oled_data = 16'b0100110001010101;
				18'b001000100110010011: oled_data = 16'b0101110100110111;
				18'b001000101000010011: oled_data = 16'b1011110100010111;
				18'b001000101010010011: oled_data = 16'b1110010010110110;
				18'b001000101100010011: oled_data = 16'b1101010001110100;
				18'b001000101110010011: oled_data = 16'b1110010011010110;
				18'b001000110000010011: oled_data = 16'b1101110011010101;
				18'b001000110010010011: oled_data = 16'b1101110011010110;
				18'b001000110100010011: oled_data = 16'b1100110000010011;
				18'b001000110110010011: oled_data = 16'b1101110010110101;
				18'b001000111000010011: oled_data = 16'b1101110011010101;
				18'b001000111010010011: oled_data = 16'b1101110011010101;
				18'b001000111100010011: oled_data = 16'b1101110011010101;
				18'b001000111110010011: oled_data = 16'b1101110011010101;
				18'b001001000000010011: oled_data = 16'b1101110011010110;
				18'b001001000010010011: oled_data = 16'b1101010010010101;
				18'b001001000100010011: oled_data = 16'b1101010010010101;
				18'b001001000110010011: oled_data = 16'b1101110011010110;
				18'b001001001000010011: oled_data = 16'b1101110011010101;
				18'b001001001010010011: oled_data = 16'b1101110011010101;
				18'b001001001100010011: oled_data = 16'b1101110010110101;
				18'b001001001110010011: oled_data = 16'b1100110000110011;
				18'b001001010000010011: oled_data = 16'b1110010011010110;
				18'b001001010010010011: oled_data = 16'b1101110011010101;
				18'b001001010100010011: oled_data = 16'b1101110011010101;
				18'b001001010110010011: oled_data = 16'b1101010001110100;
				18'b001001011000010011: oled_data = 16'b1101110011010101;
				18'b001001011010010011: oled_data = 16'b1101110011010101;
				18'b001001011100010011: oled_data = 16'b1101110011010101;
				18'b001001011110010011: oled_data = 16'b1101110011010101;
				18'b001001100000010011: oled_data = 16'b1101110011010101;
				18'b001001100010010011: oled_data = 16'b1101110011010101;
				18'b001001100100010011: oled_data = 16'b1101110011010101;
				18'b001001100110010011: oled_data = 16'b1101110011010101;
				18'b001001101000010011: oled_data = 16'b1101110011010101;
				18'b001001101010010011: oled_data = 16'b1101110011010110;
				18'b001001101100010011: oled_data = 16'b1101010001110100;
				18'b001001101110010011: oled_data = 16'b1101110010010101;
				18'b001001110000010011: oled_data = 16'b1101110011010110;
				18'b001001110010010011: oled_data = 16'b1110010011010110;
				18'b001001110100010011: oled_data = 16'b1101010010010100;
				18'b001001110110010011: oled_data = 16'b1100110001110100;
				18'b001001111000010011: oled_data = 16'b1101110011010110;
				18'b001001111010010011: oled_data = 16'b1101110011010101;
				18'b001001111100010011: oled_data = 16'b1101110011010110;
				18'b001001111110010011: oled_data = 16'b1011101110110001;
				18'b001010000000010011: oled_data = 16'b1101110010110101;
				18'b001010000010010011: oled_data = 16'b1101110011010110;
				18'b001010000100010011: oled_data = 16'b1101110011010110;
				18'b001010000110010011: oled_data = 16'b1101010001110100;
				18'b001010001000010011: oled_data = 16'b1101110010110101;
				18'b001010001010010011: oled_data = 16'b1101110011110101;
				18'b001010001100010011: oled_data = 16'b1110010100010100;
				18'b001010001110010011: oled_data = 16'b1101110001010001;
				18'b001010010000010011: oled_data = 16'b1011101010001010;
				18'b001010010010010011: oled_data = 16'b1011001000101001;
				18'b001010010100010011: oled_data = 16'b1011001001001001;
				18'b001010010110010011: oled_data = 16'b1011001001001001;
				18'b001010011000010011: oled_data = 16'b1011001001001001;
				18'b001010011010010011: oled_data = 16'b1011001000101001;
				18'b001010011100010011: oled_data = 16'b1011001001001001;
				18'b001010011110010011: oled_data = 16'b1011001000101001;
				18'b001010100000010011: oled_data = 16'b1011001000101001;
				18'b001010100010010011: oled_data = 16'b1011001000101001;
				18'b001010100100010011: oled_data = 16'b1011001000101000;
				18'b001010100110010011: oled_data = 16'b1011001000001000;
				18'b001000011000010100: oled_data = 16'b0111010111111010;
				18'b001000011010010100: oled_data = 16'b0100110010110110;
				18'b001000011100010100: oled_data = 16'b0100110001110110;
				18'b001000011110010100: oled_data = 16'b0100110001010110;
				18'b001000100000010100: oled_data = 16'b0100110001010110;
				18'b001000100010010100: oled_data = 16'b0100110001010101;
				18'b001000100100010100: oled_data = 16'b0100010001010101;
				18'b001000100110010100: oled_data = 16'b0110010100110111;
				18'b001000101000010100: oled_data = 16'b1100110010110110;
				18'b001000101010010100: oled_data = 16'b1101110010010101;
				18'b001000101100010100: oled_data = 16'b1101010010010101;
				18'b001000101110010100: oled_data = 16'b1110010011010110;
				18'b001000110000010100: oled_data = 16'b1101110011010110;
				18'b001000110010010100: oled_data = 16'b1101010010010100;
				18'b001000110100010100: oled_data = 16'b1101010001010100;
				18'b001000110110010100: oled_data = 16'b1110010011010110;
				18'b001000111000010100: oled_data = 16'b1101110011010101;
				18'b001000111010010100: oled_data = 16'b1101110011010101;
				18'b001000111100010100: oled_data = 16'b1101110011010101;
				18'b001000111110010100: oled_data = 16'b1101110011010101;
				18'b001001000000010100: oled_data = 16'b1101110011010110;
				18'b001001000010010100: oled_data = 16'b1101010010010100;
				18'b001001000100010100: oled_data = 16'b1101110010110101;
				18'b001001000110010100: oled_data = 16'b1101110011010101;
				18'b001001001000010100: oled_data = 16'b1101110011010101;
				18'b001001001010010100: oled_data = 16'b1101110011010110;
				18'b001001001100010100: oled_data = 16'b1101010010010100;
				18'b001001001110010100: oled_data = 16'b1101010001010100;
				18'b001001010000010100: oled_data = 16'b1101110011010110;
				18'b001001010010010100: oled_data = 16'b1101110011010101;
				18'b001001010100010100: oled_data = 16'b1101110010110101;
				18'b001001010110010100: oled_data = 16'b1100110000110011;
				18'b001001011000010100: oled_data = 16'b1101110011010110;
				18'b001001011010010100: oled_data = 16'b1101110011010101;
				18'b001001011100010100: oled_data = 16'b1101110011010101;
				18'b001001011110010100: oled_data = 16'b1101110011010101;
				18'b001001100000010100: oled_data = 16'b1101110011010101;
				18'b001001100010010100: oled_data = 16'b1101110011010101;
				18'b001001100100010100: oled_data = 16'b1101110011010101;
				18'b001001100110010100: oled_data = 16'b1101110011010101;
				18'b001001101000010100: oled_data = 16'b1101110011010101;
				18'b001001101010010100: oled_data = 16'b1101110011010110;
				18'b001001101100010100: oled_data = 16'b1100110001010011;
				18'b001001101110010100: oled_data = 16'b1101010010010101;
				18'b001001110000010100: oled_data = 16'b1101110011010101;
				18'b001001110010010100: oled_data = 16'b1101110010110101;
				18'b001001110100010100: oled_data = 16'b1101010010110101;
				18'b001001110110010100: oled_data = 16'b1100110010010100;
				18'b001001111000010100: oled_data = 16'b1101110011010110;
				18'b001001111010010100: oled_data = 16'b1101110011010101;
				18'b001001111100010100: oled_data = 16'b1101110010110101;
				18'b001001111110010100: oled_data = 16'b1011001110010001;
				18'b001010000000010100: oled_data = 16'b1101010010010100;
				18'b001010000010010100: oled_data = 16'b1101110011010110;
				18'b001010000100010100: oled_data = 16'b1101110011010110;
				18'b001010000110010100: oled_data = 16'b1101010010010100;
				18'b001010001000010100: oled_data = 16'b1101010001010011;
				18'b001010001010010100: oled_data = 16'b1110010011010100;
				18'b001010001100010100: oled_data = 16'b1110010010110011;
				18'b001010001110010100: oled_data = 16'b1011101010101011;
				18'b001010010000010100: oled_data = 16'b1011001001001001;
				18'b001010010010010100: oled_data = 16'b1011101001001001;
				18'b001010010100010100: oled_data = 16'b1011001001001001;
				18'b001010010110010100: oled_data = 16'b1011001001001001;
				18'b001010011000010100: oled_data = 16'b1011001001001001;
				18'b001010011010010100: oled_data = 16'b1011001000101001;
				18'b001010011100010100: oled_data = 16'b1011001001001001;
				18'b001010011110010100: oled_data = 16'b1011001000101001;
				18'b001010100000010100: oled_data = 16'b1010101000001000;
				18'b001010100010010100: oled_data = 16'b1011001000101001;
				18'b001010100100010100: oled_data = 16'b1011001000101000;
				18'b001010100110010100: oled_data = 16'b1011001000001000;
				18'b001000011000010101: oled_data = 16'b0111010110111001;
				18'b001000011010010101: oled_data = 16'b0100110010110101;
				18'b001000011100010101: oled_data = 16'b0100010001010100;
				18'b001000011110010101: oled_data = 16'b0100010001010101;
				18'b001000100000010101: oled_data = 16'b0100110001010110;
				18'b001000100010010101: oled_data = 16'b0100010001010110;
				18'b001000100100010101: oled_data = 16'b0100110010010110;
				18'b001000100110010101: oled_data = 16'b1000010100010111;
				18'b001000101000010101: oled_data = 16'b1101010010010101;
				18'b001000101010010101: oled_data = 16'b1101010001110100;
				18'b001000101100010101: oled_data = 16'b1101110011010101;
				18'b001000101110010101: oled_data = 16'b1101110011010101;
				18'b001000110000010101: oled_data = 16'b1101110011010101;
				18'b001000110010010101: oled_data = 16'b1100110001010011;
				18'b001000110100010101: oled_data = 16'b1101010010010101;
				18'b001000110110010101: oled_data = 16'b1110010011110110;
				18'b001000111000010101: oled_data = 16'b1101110011010101;
				18'b001000111010010101: oled_data = 16'b1101110011010101;
				18'b001000111100010101: oled_data = 16'b1101110011010101;
				18'b001000111110010101: oled_data = 16'b1101110011010101;
				18'b001001000000010101: oled_data = 16'b1101110011010101;
				18'b001001000010010101: oled_data = 16'b1101010001110100;
				18'b001001000100010101: oled_data = 16'b1101110011010101;
				18'b001001000110010101: oled_data = 16'b1101110011010101;
				18'b001001001000010101: oled_data = 16'b1101110011010101;
				18'b001001001010010101: oled_data = 16'b1110010011110110;
				18'b001001001100010101: oled_data = 16'b1100110001110100;
				18'b001001001110010101: oled_data = 16'b1101010010010100;
				18'b001001010000010101: oled_data = 16'b1101110011010110;
				18'b001001010010010101: oled_data = 16'b1101110011010110;
				18'b001001010100010101: oled_data = 16'b1101010010110101;
				18'b001001010110010101: oled_data = 16'b1100110001010011;
				18'b001001011000010101: oled_data = 16'b1101110011010110;
				18'b001001011010010101: oled_data = 16'b1101110011010101;
				18'b001001011100010101: oled_data = 16'b1101110011010101;
				18'b001001011110010101: oled_data = 16'b1101110011010101;
				18'b001001100000010101: oled_data = 16'b1101110011010101;
				18'b001001100010010101: oled_data = 16'b1101110011010101;
				18'b001001100100010101: oled_data = 16'b1101110011010101;
				18'b001001100110010101: oled_data = 16'b1101110011010101;
				18'b001001101000010101: oled_data = 16'b1101110010110101;
				18'b001001101010010101: oled_data = 16'b1101110011010101;
				18'b001001101100010101: oled_data = 16'b1101010001110100;
				18'b001001101110010101: oled_data = 16'b1101110010110101;
				18'b001001110000010101: oled_data = 16'b1101010010010101;
				18'b001001110010010101: oled_data = 16'b1101010010010101;
				18'b001001110100010101: oled_data = 16'b1101010011010101;
				18'b001001110110010101: oled_data = 16'b1101010010110100;
				18'b001001111000010101: oled_data = 16'b1110010011010101;
				18'b001001111010010101: oled_data = 16'b1101110011010110;
				18'b001001111100010101: oled_data = 16'b1101110010010101;
				18'b001001111110010101: oled_data = 16'b1011001101010000;
				18'b001010000000010101: oled_data = 16'b1101010001110100;
				18'b001010000010010101: oled_data = 16'b1101110011010110;
				18'b001010000100010101: oled_data = 16'b1101110011010110;
				18'b001010000110010101: oled_data = 16'b1101010001110100;
				18'b001010001000010101: oled_data = 16'b1101010010010011;
				18'b001010001010010101: oled_data = 16'b1110110011110100;
				18'b001010001100010101: oled_data = 16'b1100001100101101;
				18'b001010001110010101: oled_data = 16'b1011001000101001;
				18'b001010010000010101: oled_data = 16'b1011101001001001;
				18'b001010010010010101: oled_data = 16'b1011101000101001;
				18'b001010010100010101: oled_data = 16'b1011001001001001;
				18'b001010010110010101: oled_data = 16'b1011001001001001;
				18'b001010011000010101: oled_data = 16'b1011001001001001;
				18'b001010011010010101: oled_data = 16'b1011001001001001;
				18'b001010011100010101: oled_data = 16'b1011001000101001;
				18'b001010011110010101: oled_data = 16'b1010001000001000;
				18'b001010100000010101: oled_data = 16'b1010101000001000;
				18'b001010100010010101: oled_data = 16'b1011001000101001;
				18'b001010100100010101: oled_data = 16'b1011001000101000;
				18'b001010100110010101: oled_data = 16'b1011001000001000;
				18'b001000011000010110: oled_data = 16'b1010010011110100;
				18'b001000011010010110: oled_data = 16'b0111010001110100;
				18'b001000011100010110: oled_data = 16'b0100110001110101;
				18'b001000011110010110: oled_data = 16'b0100010001110110;
				18'b001000100000010110: oled_data = 16'b0100010001110101;
				18'b001000100010010110: oled_data = 16'b0100010001110101;
				18'b001000100100010110: oled_data = 16'b0110010101011000;
				18'b001000100110010110: oled_data = 16'b1010110010110110;
				18'b001000101000010110: oled_data = 16'b1101010010010101;
				18'b001000101010010110: oled_data = 16'b1101010010010101;
				18'b001000101100010110: oled_data = 16'b1101110011010101;
				18'b001000101110010110: oled_data = 16'b1101110011010110;
				18'b001000110000010110: oled_data = 16'b1101110010010101;
				18'b001000110010010110: oled_data = 16'b1101010001110100;
				18'b001000110100010110: oled_data = 16'b1101010010110101;
				18'b001000110110010110: oled_data = 16'b1101110011110110;
				18'b001000111000010110: oled_data = 16'b1101110011010101;
				18'b001000111010010110: oled_data = 16'b1101110011010101;
				18'b001000111100010110: oled_data = 16'b1101110011010101;
				18'b001000111110010110: oled_data = 16'b1101110011010101;
				18'b001001000000010110: oled_data = 16'b1101110010110101;
				18'b001001000010010110: oled_data = 16'b1101010001110100;
				18'b001001000100010110: oled_data = 16'b1101110011010110;
				18'b001001000110010110: oled_data = 16'b1101110011010101;
				18'b001001001000010110: oled_data = 16'b1101110011010101;
				18'b001001001010010110: oled_data = 16'b1101110011010110;
				18'b001001001100010110: oled_data = 16'b1100110001110100;
				18'b001001001110010110: oled_data = 16'b1101110010110101;
				18'b001001010000010110: oled_data = 16'b1101110011010101;
				18'b001001010010010110: oled_data = 16'b1101110011010110;
				18'b001001010100010110: oled_data = 16'b1101010010010100;
				18'b001001010110010110: oled_data = 16'b1100110010010100;
				18'b001001011000010110: oled_data = 16'b1101110011010110;
				18'b001001011010010110: oled_data = 16'b1101110011010101;
				18'b001001011100010110: oled_data = 16'b1101110011010101;
				18'b001001011110010110: oled_data = 16'b1101110011010101;
				18'b001001100000010110: oled_data = 16'b1101110011010101;
				18'b001001100010010110: oled_data = 16'b1101110011010101;
				18'b001001100100010110: oled_data = 16'b1101110011010101;
				18'b001001100110010110: oled_data = 16'b1101110011010110;
				18'b001001101000010110: oled_data = 16'b1101010010010100;
				18'b001001101010010110: oled_data = 16'b1101110011010101;
				18'b001001101100010110: oled_data = 16'b1101010001110100;
				18'b001001101110010110: oled_data = 16'b1101010010010100;
				18'b001001110000010110: oled_data = 16'b1101110010110101;
				18'b001001110010010110: oled_data = 16'b1011110000010010;
				18'b001001110100010110: oled_data = 16'b0111001010101011;
				18'b001001110110010110: oled_data = 16'b1100110010110011;
				18'b001001111000010110: oled_data = 16'b1110010011010101;
				18'b001001111010010110: oled_data = 16'b1101110011010110;
				18'b001001111100010110: oled_data = 16'b1100110001010100;
				18'b001001111110010110: oled_data = 16'b1010101100101111;
				18'b001010000000010110: oled_data = 16'b1100110001010100;
				18'b001010000010010110: oled_data = 16'b1101110011110110;
				18'b001010000100010110: oled_data = 16'b1101110011010101;
				18'b001010000110010110: oled_data = 16'b1101010001110011;
				18'b001010001000010110: oled_data = 16'b1110110100010100;
				18'b001010001010010110: oled_data = 16'b1101001111101111;
				18'b001010001100010110: oled_data = 16'b1011001001001001;
				18'b001010001110010110: oled_data = 16'b1011101001001001;
				18'b001010010000010110: oled_data = 16'b1011101001001001;
				18'b001010010010010110: oled_data = 16'b1011101001001001;
				18'b001010010100010110: oled_data = 16'b1011001001001001;
				18'b001010010110010110: oled_data = 16'b1011001001001001;
				18'b001010011000010110: oled_data = 16'b1011001001001001;
				18'b001010011010010110: oled_data = 16'b1010101000101000;
				18'b001010011100010110: oled_data = 16'b1010001000001000;
				18'b001010011110010110: oled_data = 16'b1011001000101001;
				18'b001010100000010110: oled_data = 16'b1011001000101001;
				18'b001010100010010110: oled_data = 16'b1011001000101001;
				18'b001010100100010110: oled_data = 16'b1011001000101000;
				18'b001010100110010110: oled_data = 16'b1011001000001000;
				18'b001000011000010111: oled_data = 16'b1101011001001111;
				18'b001000011010010111: oled_data = 16'b1010110111001110;
				18'b001000011100010111: oled_data = 16'b1001010110110011;
				18'b001000011110010111: oled_data = 16'b0111010110010111;
				18'b001000100000010111: oled_data = 16'b0110010101111000;
				18'b001000100010010111: oled_data = 16'b0110010110111001;
				18'b001000100100010111: oled_data = 16'b1000010110011000;
				18'b001000100110010111: oled_data = 16'b1100110001010101;
				18'b001000101000010111: oled_data = 16'b1101010001110100;
				18'b001000101010010111: oled_data = 16'b1101110010110101;
				18'b001000101100010111: oled_data = 16'b1101110011010101;
				18'b001000101110010111: oled_data = 16'b1101110011010101;
				18'b001000110000010111: oled_data = 16'b1101010001110100;
				18'b001000110010010111: oled_data = 16'b1101010001110100;
				18'b001000110100010111: oled_data = 16'b1101110010110101;
				18'b001000110110010111: oled_data = 16'b1101110011010101;
				18'b001000111000010111: oled_data = 16'b1101110011010101;
				18'b001000111010010111: oled_data = 16'b1101110011010101;
				18'b001000111100010111: oled_data = 16'b1101110011010101;
				18'b001000111110010111: oled_data = 16'b1101110011010110;
				18'b001001000000010111: oled_data = 16'b1101010010010101;
				18'b001001000010010111: oled_data = 16'b1101110010010101;
				18'b001001000100010111: oled_data = 16'b1101110011010110;
				18'b001001000110010111: oled_data = 16'b1101110011010101;
				18'b001001001000010111: oled_data = 16'b1101110011010110;
				18'b001001001010010111: oled_data = 16'b1101110011010101;
				18'b001001001100010111: oled_data = 16'b1100110011010100;
				18'b001001001110010111: oled_data = 16'b1101110011010101;
				18'b001001010000010111: oled_data = 16'b1101110011010101;
				18'b001001010010010111: oled_data = 16'b1110010011010110;
				18'b001001010100010111: oled_data = 16'b1100110010010100;
				18'b001001010110010111: oled_data = 16'b1100110010110101;
				18'b001001011000010111: oled_data = 16'b1101110011010110;
				18'b001001011010010111: oled_data = 16'b1110010011010101;
				18'b001001011100010111: oled_data = 16'b1110010011010101;
				18'b001001011110010111: oled_data = 16'b1101110011010101;
				18'b001001100000010111: oled_data = 16'b1101110011010101;
				18'b001001100010010111: oled_data = 16'b1101110011010101;
				18'b001001100100010111: oled_data = 16'b1101110011010101;
				18'b001001100110010111: oled_data = 16'b1101110011010101;
				18'b001001101000010111: oled_data = 16'b1101010010010101;
				18'b001001101010010111: oled_data = 16'b1101110011010101;
				18'b001001101100010111: oled_data = 16'b1100010000110011;
				18'b001001101110010111: oled_data = 16'b1100110001110100;
				18'b001001110000010111: oled_data = 16'b1110010100010110;
				18'b001001110010010111: oled_data = 16'b1000101011101101;
				18'b001001110100010111: oled_data = 16'b0111001100101101;
				18'b001001110110010111: oled_data = 16'b1101010100110110;
				18'b001001111000010111: oled_data = 16'b1101110011010101;
				18'b001001111010010111: oled_data = 16'b1101110011110110;
				18'b001001111100010111: oled_data = 16'b1100001111110010;
				18'b001001111110010111: oled_data = 16'b1011001101010000;
				18'b001010000000010111: oled_data = 16'b1100110001010011;
				18'b001010000010010111: oled_data = 16'b1101110011110110;
				18'b001010000100010111: oled_data = 16'b1101010010010011;
				18'b001010000110010111: oled_data = 16'b1110010011110100;
				18'b001010001000010111: oled_data = 16'b1110010010110010;
				18'b001010001010010111: oled_data = 16'b1011101010001010;
				18'b001010001100010111: oled_data = 16'b1011001000101001;
				18'b001010001110010111: oled_data = 16'b1011001001001001;
				18'b001010010000010111: oled_data = 16'b1011001001001001;
				18'b001010010010010111: oled_data = 16'b1011001001001001;
				18'b001010010100010111: oled_data = 16'b1011001001001001;
				18'b001010010110010111: oled_data = 16'b1011001001001001;
				18'b001010011000010111: oled_data = 16'b1011001000101001;
				18'b001010011010010111: oled_data = 16'b1010001000001000;
				18'b001010011100010111: oled_data = 16'b1011001001001001;
				18'b001010011110010111: oled_data = 16'b1011001000101001;
				18'b001010100000010111: oled_data = 16'b1011001000101001;
				18'b001010100010010111: oled_data = 16'b1011001000101001;
				18'b001010100100010111: oled_data = 16'b1011001000101000;
				18'b001010100110010111: oled_data = 16'b1011001000001000;
				18'b001000011000011000: oled_data = 16'b1111011100110110;
				18'b001000011010011000: oled_data = 16'b1110011001110000;
				18'b001000011100011000: oled_data = 16'b1011110100101010;
				18'b001000011110011000: oled_data = 16'b1011010101101010;
				18'b001000100000011000: oled_data = 16'b1011011000010001;
				18'b001000100010011000: oled_data = 16'b1010010111110010;
				18'b001000100100011000: oled_data = 16'b1010010001010010;
				18'b001000100110011000: oled_data = 16'b1101110001110101;
				18'b001000101000011000: oled_data = 16'b1100110001110100;
				18'b001000101010011000: oled_data = 16'b1101110011010110;
				18'b001000101100011000: oled_data = 16'b1101110011010110;
				18'b001000101110011000: oled_data = 16'b1101010010010101;
				18'b001000110000011000: oled_data = 16'b1101010010010100;
				18'b001000110010011000: oled_data = 16'b1101010001110100;
				18'b001000110100011000: oled_data = 16'b1101110011010101;
				18'b001000110110011000: oled_data = 16'b1101110011010101;
				18'b001000111000011000: oled_data = 16'b1101110011010101;
				18'b001000111010011000: oled_data = 16'b1101110011010101;
				18'b001000111100011000: oled_data = 16'b1101110011010101;
				18'b001000111110011000: oled_data = 16'b1101110011010110;
				18'b001001000000011000: oled_data = 16'b1101010001110100;
				18'b001001000010011000: oled_data = 16'b1101110010110101;
				18'b001001000100011000: oled_data = 16'b1101110011010101;
				18'b001001000110011000: oled_data = 16'b1101110011010101;
				18'b001001001000011000: oled_data = 16'b1101110011010110;
				18'b001001001010011000: oled_data = 16'b1101010010110100;
				18'b001001001100011000: oled_data = 16'b1101010101110101;
				18'b001001001110011000: oled_data = 16'b1101110011010101;
				18'b001001010000011000: oled_data = 16'b1101110011010101;
				18'b001001010010011000: oled_data = 16'b1101110010110101;
				18'b001001010100011000: oled_data = 16'b1101010100010110;
				18'b001001010110011000: oled_data = 16'b1101010011110101;
				18'b001001011000011000: oled_data = 16'b1101110011010101;
				18'b001001011010011000: oled_data = 16'b1110010011010101;
				18'b001001011100011000: oled_data = 16'b1110010011010101;
				18'b001001011110011000: oled_data = 16'b1101110011010101;
				18'b001001100000011000: oled_data = 16'b1101110011010101;
				18'b001001100010011000: oled_data = 16'b1101110011010101;
				18'b001001100100011000: oled_data = 16'b1101110011010101;
				18'b001001100110011000: oled_data = 16'b1101110011010101;
				18'b001001101000011000: oled_data = 16'b1101010001110100;
				18'b001001101010011000: oled_data = 16'b1101010001110100;
				18'b001001101100011000: oled_data = 16'b1100010001110011;
				18'b001001101110011000: oled_data = 16'b1101110011110110;
				18'b001001110000011000: oled_data = 16'b1101110010110101;
				18'b001001110010011000: oled_data = 16'b0110000111101001;
				18'b001001110100011000: oled_data = 16'b1010110011110100;
				18'b001001110110011000: oled_data = 16'b1101110101010110;
				18'b001001111000011000: oled_data = 16'b1101110011010101;
				18'b001001111010011000: oled_data = 16'b1101110011010101;
				18'b001001111100011000: oled_data = 16'b1011101110010001;
				18'b001001111110011000: oled_data = 16'b1011001101110001;
				18'b001010000000011000: oled_data = 16'b1100110000110011;
				18'b001010000010011000: oled_data = 16'b1101110010110101;
				18'b001010000100011000: oled_data = 16'b1101010010010011;
				18'b001010000110011000: oled_data = 16'b1110110100010100;
				18'b001010001000011000: oled_data = 16'b1100101101101101;
				18'b001010001010011000: oled_data = 16'b1011001000101001;
				18'b001010001100011000: oled_data = 16'b1011001001001001;
				18'b001010001110011000: oled_data = 16'b1011001001001001;
				18'b001010010000011000: oled_data = 16'b1011001001001001;
				18'b001010010010011000: oled_data = 16'b1011001001001001;
				18'b001010010100011000: oled_data = 16'b1011001001001001;
				18'b001010010110011000: oled_data = 16'b1011001000101001;
				18'b001010011000011000: oled_data = 16'b1010101000001000;
				18'b001010011010011000: oled_data = 16'b1011001000101001;
				18'b001010011100011000: oled_data = 16'b1011001001001001;
				18'b001010011110011000: oled_data = 16'b1011001000101001;
				18'b001010100000011000: oled_data = 16'b1011001000101001;
				18'b001010100010011000: oled_data = 16'b1011001000101001;
				18'b001010100100011000: oled_data = 16'b1011001000101000;
				18'b001010100110011000: oled_data = 16'b1010101000001000;
				18'b001000011000011001: oled_data = 16'b1101011000001111;
				18'b001000011010011001: oled_data = 16'b1101010111101111;
				18'b001000011100011001: oled_data = 16'b1011010100001010;
				18'b001000011110011001: oled_data = 16'b1010110010100111;
				18'b001000100000011001: oled_data = 16'b1100010110001001;
				18'b001000100010011001: oled_data = 16'b1101011001001011;
				18'b001000100100011001: oled_data = 16'b1100110010010000;
				18'b001000100110011001: oled_data = 16'b1101110010010101;
				18'b001000101000011001: oled_data = 16'b1101010010010101;
				18'b001000101010011001: oled_data = 16'b1101110011010110;
				18'b001000101100011001: oled_data = 16'b1101110011010110;
				18'b001000101110011001: oled_data = 16'b1101010001110100;
				18'b001000110000011001: oled_data = 16'b1101110011010101;
				18'b001000110010011001: oled_data = 16'b1101010001110100;
				18'b001000110100011001: oled_data = 16'b1110010011010110;
				18'b001000110110011001: oled_data = 16'b1101110011010101;
				18'b001000111000011001: oled_data = 16'b1101110011010101;
				18'b001000111010011001: oled_data = 16'b1101110011010101;
				18'b001000111100011001: oled_data = 16'b1101110011010101;
				18'b001000111110011001: oled_data = 16'b1101110011010101;
				18'b001001000000011001: oled_data = 16'b1101010001110100;
				18'b001001000010011001: oled_data = 16'b1101110011010101;
				18'b001001000100011001: oled_data = 16'b1101110011010101;
				18'b001001000110011001: oled_data = 16'b1101110011010101;
				18'b001001001000011001: oled_data = 16'b1101110010110101;
				18'b001001001010011001: oled_data = 16'b1101010100010101;
				18'b001001001100011001: oled_data = 16'b1101111000111000;
				18'b001001001110011001: oled_data = 16'b1101110011010101;
				18'b001001010000011001: oled_data = 16'b1110010011010110;
				18'b001001010010011001: oled_data = 16'b1101110010110101;
				18'b001001010100011001: oled_data = 16'b1101110111011000;
				18'b001001010110011001: oled_data = 16'b1101110011110110;
				18'b001001011000011001: oled_data = 16'b1101110011010101;
				18'b001001011010011001: oled_data = 16'b1101110011010101;
				18'b001001011100011001: oled_data = 16'b1101110011010101;
				18'b001001011110011001: oled_data = 16'b1101110011010101;
				18'b001001100000011001: oled_data = 16'b1101110011010101;
				18'b001001100010011001: oled_data = 16'b1101110011010101;
				18'b001001100100011001: oled_data = 16'b1101110011010101;
				18'b001001100110011001: oled_data = 16'b1101110010110101;
				18'b001001101000011001: oled_data = 16'b1101010001110100;
				18'b001001101010011001: oled_data = 16'b1101010011110101;
				18'b001001101100011001: oled_data = 16'b1101010100110101;
				18'b001001101110011001: oled_data = 16'b1110010011010110;
				18'b001001110000011001: oled_data = 16'b1011001111010001;
				18'b001001110010011001: oled_data = 16'b0101101000001001;
				18'b001001110100011001: oled_data = 16'b1101011001011001;
				18'b001001110110011001: oled_data = 16'b1101010100110110;
				18'b001001111000011001: oled_data = 16'b1110010011010110;
				18'b001001111010011001: oled_data = 16'b1101010001010100;
				18'b001001111100011001: oled_data = 16'b1011001101010000;
				18'b001001111110011001: oled_data = 16'b1011001101110001;
				18'b001010000000011001: oled_data = 16'b1100110000110011;
				18'b001010000010011001: oled_data = 16'b1101010010010100;
				18'b001010000100011001: oled_data = 16'b1110010100010100;
				18'b001010000110011001: oled_data = 16'b1101110001110001;
				18'b001010001000011001: oled_data = 16'b1011101001101010;
				18'b001010001010011001: oled_data = 16'b1011001001001001;
				18'b001010001100011001: oled_data = 16'b1011001001001001;
				18'b001010001110011001: oled_data = 16'b1011001001001001;
				18'b001010010000011001: oled_data = 16'b1011001001001001;
				18'b001010010010011001: oled_data = 16'b1011001001001001;
				18'b001010010100011001: oled_data = 16'b1011001000101001;
				18'b001010010110011001: oled_data = 16'b1010101000001000;
				18'b001010011000011001: oled_data = 16'b1011001000101001;
				18'b001010011010011001: oled_data = 16'b1011001001001001;
				18'b001010011100011001: oled_data = 16'b1011001000101001;
				18'b001010011110011001: oled_data = 16'b1011001000101001;
				18'b001010100000011001: oled_data = 16'b1011001000101001;
				18'b001010100010011001: oled_data = 16'b1011001000101000;
				18'b001010100100011001: oled_data = 16'b1011001000101000;
				18'b001010100110011001: oled_data = 16'b1010101000101000;
				18'b001000011000011010: oled_data = 16'b1010010010101000;
				18'b001000011010011010: oled_data = 16'b1010010010001000;
				18'b001000011100011010: oled_data = 16'b1010110010101000;
				18'b001000011110011010: oled_data = 16'b1010110010101000;
				18'b001000100000011010: oled_data = 16'b1010110011101000;
				18'b001000100010011010: oled_data = 16'b1100111000001011;
				18'b001000100100011010: oled_data = 16'b1101010100010001;
				18'b001000100110011010: oled_data = 16'b1101010001110100;
				18'b001000101000011010: oled_data = 16'b1101110011010101;
				18'b001000101010011010: oled_data = 16'b1101110011010110;
				18'b001000101100011010: oled_data = 16'b1101110011010101;
				18'b001000101110011010: oled_data = 16'b1101010010010100;
				18'b001000110000011010: oled_data = 16'b1110010011010110;
				18'b001000110010011010: oled_data = 16'b1101010010010100;
				18'b001000110100011010: oled_data = 16'b1110010011110110;
				18'b001000110110011010: oled_data = 16'b1101110011010101;
				18'b001000111000011010: oled_data = 16'b1101110011010101;
				18'b001000111010011010: oled_data = 16'b1101110011010101;
				18'b001000111100011010: oled_data = 16'b1101110011010101;
				18'b001000111110011010: oled_data = 16'b1101110010110101;
				18'b001001000000011010: oled_data = 16'b1101010001110100;
				18'b001001000010011010: oled_data = 16'b1101110011010110;
				18'b001001000100011010: oled_data = 16'b1101110011010101;
				18'b001001000110011010: oled_data = 16'b1101110011010101;
				18'b001001001000011010: oled_data = 16'b1101110010010101;
				18'b001001001010011010: oled_data = 16'b1101110110110111;
				18'b001001001100011010: oled_data = 16'b1110011001011000;
				18'b001001001110011010: oled_data = 16'b1101110011010101;
				18'b001001010000011010: oled_data = 16'b1101110011010101;
				18'b001001010010011010: oled_data = 16'b1101010011010101;
				18'b001001010100011010: oled_data = 16'b1101111001011001;
				18'b001001010110011010: oled_data = 16'b1101110011110110;
				18'b001001011000011010: oled_data = 16'b1101110011010110;
				18'b001001011010011010: oled_data = 16'b1101110010110101;
				18'b001001011100011010: oled_data = 16'b1101110010110101;
				18'b001001011110011010: oled_data = 16'b1101110011010101;
				18'b001001100000011010: oled_data = 16'b1101110011010101;
				18'b001001100010011010: oled_data = 16'b1101110011010101;
				18'b001001100100011010: oled_data = 16'b1101110011010110;
				18'b001001100110011010: oled_data = 16'b1101010010010101;
				18'b001001101000011010: oled_data = 16'b1101110010010101;
				18'b001001101010011010: oled_data = 16'b1101010100110110;
				18'b001001101100011010: oled_data = 16'b1100110101010101;
				18'b001001101110011010: oled_data = 16'b1110010011010101;
				18'b001001110000011010: oled_data = 16'b1000101010001100;
				18'b001001110010011010: oled_data = 16'b0111101101001110;
				18'b001001110100011010: oled_data = 16'b1110111100011100;
				18'b001001110110011010: oled_data = 16'b1101010100010110;
				18'b001001111000011010: oled_data = 16'b1101110011010110;
				18'b001001111010011010: oled_data = 16'b1100010000110011;
				18'b001001111100011010: oled_data = 16'b1011001101110001;
				18'b001001111110011010: oled_data = 16'b1011101101110001;
				18'b001010000000011010: oled_data = 16'b1100110000010010;
				18'b001010000010011010: oled_data = 16'b1101110010110011;
				18'b001010000100011010: oled_data = 16'b1110110100010100;
				18'b001010000110011010: oled_data = 16'b1100101100101101;
				18'b001010001000011010: oled_data = 16'b1011001001001001;
				18'b001010001010011010: oled_data = 16'b1011001001001001;
				18'b001010001100011010: oled_data = 16'b1011001001001001;
				18'b001010001110011010: oled_data = 16'b1011001001001001;
				18'b001010010000011010: oled_data = 16'b1011001001001001;
				18'b001010010010011010: oled_data = 16'b1011001001001001;
				18'b001010010100011010: oled_data = 16'b1010101000001000;
				18'b001010010110011010: oled_data = 16'b1011001000101001;
				18'b001010011000011010: oled_data = 16'b1011001001001001;
				18'b001010011010011010: oled_data = 16'b1011001001001001;
				18'b001010011100011010: oled_data = 16'b1011001000101001;
				18'b001010011110011010: oled_data = 16'b1011001000101001;
				18'b001010100000011010: oled_data = 16'b1011001000101001;
				18'b001010100010011010: oled_data = 16'b1011001000101000;
				18'b001010100100011010: oled_data = 16'b1011001000101000;
				18'b001010100110011010: oled_data = 16'b1010101000101000;
				18'b001000011000011011: oled_data = 16'b1010110010100111;
				18'b001000011010011011: oled_data = 16'b1010110010100111;
				18'b001000011100011011: oled_data = 16'b1010110010101000;
				18'b001000011110011011: oled_data = 16'b1010110010101000;
				18'b001000100000011011: oled_data = 16'b1010110010100111;
				18'b001000100010011011: oled_data = 16'b1100110110101010;
				18'b001000100100011011: oled_data = 16'b1101010100010001;
				18'b001000100110011011: oled_data = 16'b1101010001110100;
				18'b001000101000011011: oled_data = 16'b1101110011010101;
				18'b001000101010011011: oled_data = 16'b1101110011010110;
				18'b001000101100011011: oled_data = 16'b1101010010010101;
				18'b001000101110011011: oled_data = 16'b1101110010110101;
				18'b001000110000011011: oled_data = 16'b1101110011010101;
				18'b001000110010011011: oled_data = 16'b1101110010110101;
				18'b001000110100011011: oled_data = 16'b1110010011110110;
				18'b001000110110011011: oled_data = 16'b1101110011010101;
				18'b001000111000011011: oled_data = 16'b1101110011010101;
				18'b001000111010011011: oled_data = 16'b1101110011010101;
				18'b001000111100011011: oled_data = 16'b1101110011010101;
				18'b001000111110011011: oled_data = 16'b1101110010110101;
				18'b001001000000011011: oled_data = 16'b1101010010010100;
				18'b001001000010011011: oled_data = 16'b1101110011010110;
				18'b001001000100011011: oled_data = 16'b1101110011010101;
				18'b001001000110011011: oled_data = 16'b1110010011010101;
				18'b001001001000011011: oled_data = 16'b1101010011010101;
				18'b001001001010011011: oled_data = 16'b1110011010011010;
				18'b001001001100011011: oled_data = 16'b1101111001111000;
				18'b001001001110011011: oled_data = 16'b1101110011010101;
				18'b001001010000011011: oled_data = 16'b1110010011010110;
				18'b001001010010011011: oled_data = 16'b1101010100010110;
				18'b001001010100011011: oled_data = 16'b1110011010011010;
				18'b001001010110011011: oled_data = 16'b1101010011110101;
				18'b001001011000011011: oled_data = 16'b1110010011110110;
				18'b001001011010011011: oled_data = 16'b1101010001110100;
				18'b001001011100011011: oled_data = 16'b1101110010110101;
				18'b001001011110011011: oled_data = 16'b1101110011010101;
				18'b001001100000011011: oled_data = 16'b1101110011010101;
				18'b001001100010011011: oled_data = 16'b1101110011010101;
				18'b001001100100011011: oled_data = 16'b1101110011010110;
				18'b001001100110011011: oled_data = 16'b1101010001110100;
				18'b001001101000011011: oled_data = 16'b1101110010110101;
				18'b001001101010011011: oled_data = 16'b1101110111011000;
				18'b001001101100011011: oled_data = 16'b1101010101110110;
				18'b001001101110011011: oled_data = 16'b1100110010010011;
				18'b001001110000011011: oled_data = 16'b0101100111001000;
				18'b001001110010011011: oled_data = 16'b1011010101010100;
				18'b001001110100011011: oled_data = 16'b1110111011111011;
				18'b001001110110011011: oled_data = 16'b1101010011110101;
				18'b001001111000011011: oled_data = 16'b1101010011010101;
				18'b001001111010011011: oled_data = 16'b1101110111111000;
				18'b001001111100011011: oled_data = 16'b1011001111110001;
				18'b001001111110011011: oled_data = 16'b1011001101110001;
				18'b001010000000011011: oled_data = 16'b1011101111010001;
				18'b001010000010011011: oled_data = 16'b1110110100010100;
				18'b001010000100011011: oled_data = 16'b1110010001110001;
				18'b001010000110011011: oled_data = 16'b1011101001101010;
				18'b001010001000011011: oled_data = 16'b1011101001001001;
				18'b001010001010011011: oled_data = 16'b1100001011001100;
				18'b001010001100011011: oled_data = 16'b1011101001101010;
				18'b001010001110011011: oled_data = 16'b1011001001001001;
				18'b001010010000011011: oled_data = 16'b1011001001001001;
				18'b001010010010011011: oled_data = 16'b1011001000101000;
				18'b001010010100011011: oled_data = 16'b1010101000101001;
				18'b001010010110011011: oled_data = 16'b1011001001001001;
				18'b001010011000011011: oled_data = 16'b1011001001001001;
				18'b001010011010011011: oled_data = 16'b1011001000101001;
				18'b001010011100011011: oled_data = 16'b1011001000101001;
				18'b001010011110011011: oled_data = 16'b1011001000101001;
				18'b001010100000011011: oled_data = 16'b1011001000101001;
				18'b001010100010011011: oled_data = 16'b1011001000101000;
				18'b001010100100011011: oled_data = 16'b1011001000101000;
				18'b001010100110011011: oled_data = 16'b1010101000101000;
				18'b001000011000011100: oled_data = 16'b1010110010100111;
				18'b001000011010011100: oled_data = 16'b1010110010100111;
				18'b001000011100011100: oled_data = 16'b1010110010101000;
				18'b001000011110011100: oled_data = 16'b1010110010101000;
				18'b001000100000011100: oled_data = 16'b1010110010100111;
				18'b001000100010011100: oled_data = 16'b1100010101101010;
				18'b001000100100011100: oled_data = 16'b1101010011110010;
				18'b001000100110011100: oled_data = 16'b1101110010010101;
				18'b001000101000011100: oled_data = 16'b1101110011010110;
				18'b001000101010011100: oled_data = 16'b1101110011010101;
				18'b001000101100011100: oled_data = 16'b1101010010010100;
				18'b001000101110011100: oled_data = 16'b1101110011010101;
				18'b001000110000011100: oled_data = 16'b1101110011010101;
				18'b001000110010011100: oled_data = 16'b1101010010010100;
				18'b001000110100011100: oled_data = 16'b1110010011110110;
				18'b001000110110011100: oled_data = 16'b1101110011010101;
				18'b001000111000011100: oled_data = 16'b1101110011010101;
				18'b001000111010011100: oled_data = 16'b1101110011010101;
				18'b001000111100011100: oled_data = 16'b1101110011010110;
				18'b001000111110011100: oled_data = 16'b1101110010010101;
				18'b001001000000011100: oled_data = 16'b1101110010010101;
				18'b001001000010011100: oled_data = 16'b1101110011010110;
				18'b001001000100011100: oled_data = 16'b1101110011010101;
				18'b001001000110011100: oled_data = 16'b1101110010110101;
				18'b001001001000011100: oled_data = 16'b1101110101110111;
				18'b001001001010011100: oled_data = 16'b1110111011111011;
				18'b001001001100011100: oled_data = 16'b1101111001011000;
				18'b001001001110011100: oled_data = 16'b1101110011010101;
				18'b001001010000011100: oled_data = 16'b1101110011010110;
				18'b001001010010011100: oled_data = 16'b1101110110010111;
				18'b001001010100011100: oled_data = 16'b1101111010011010;
				18'b001001010110011100: oled_data = 16'b1101010011110101;
				18'b001001011000011100: oled_data = 16'b1101110011010101;
				18'b001001011010011100: oled_data = 16'b1101010001110100;
				18'b001001011100011100: oled_data = 16'b1101110011010101;
				18'b001001011110011100: oled_data = 16'b1101110011010101;
				18'b001001100000011100: oled_data = 16'b1101110011010101;
				18'b001001100010011100: oled_data = 16'b1101110011010101;
				18'b001001100100011100: oled_data = 16'b1101110010110101;
				18'b001001100110011100: oled_data = 16'b1101010001110100;
				18'b001001101000011100: oled_data = 16'b1101110011010101;
				18'b001001101010011100: oled_data = 16'b1101111000111001;
				18'b001001101100011100: oled_data = 16'b1101010101110110;
				18'b001001101110011100: oled_data = 16'b1010001110001111;
				18'b001001110000011100: oled_data = 16'b0100100111101000;
				18'b001001110010011100: oled_data = 16'b1101111011011010;
				18'b001001110100011100: oled_data = 16'b1101111010111010;
				18'b001001110110011100: oled_data = 16'b1101010011010101;
				18'b001001111000011100: oled_data = 16'b1101110110010111;
				18'b001001111010011100: oled_data = 16'b1110111100111011;
				18'b001001111100011100: oled_data = 16'b1100010011010100;
				18'b001001111110011100: oled_data = 16'b1011001100101111;
				18'b001010000000011100: oled_data = 16'b1100110000110001;
				18'b001010000010011100: oled_data = 16'b1110110100010100;
				18'b001010000100011100: oled_data = 16'b1100101101101101;
				18'b001010000110011100: oled_data = 16'b1011001000101001;
				18'b001010001000011100: oled_data = 16'b1011101010001010;
				18'b001010001010011100: oled_data = 16'b1101001110001110;
				18'b001010001100011100: oled_data = 16'b1011001001001010;
				18'b001010001110011100: oled_data = 16'b1011101001001001;
				18'b001010010000011100: oled_data = 16'b1011001001001001;
				18'b001010010010011100: oled_data = 16'b1010101000001000;
				18'b001010010100011100: oled_data = 16'b1011101001001001;
				18'b001010010110011100: oled_data = 16'b1011001001001001;
				18'b001010011000011100: oled_data = 16'b1010000111101000;
				18'b001010011010011100: oled_data = 16'b1010000111000111;
				18'b001010011100011100: oled_data = 16'b1011001001001001;
				18'b001010011110011100: oled_data = 16'b1011001000101000;
				18'b001010100000011100: oled_data = 16'b1011001000101001;
				18'b001010100010011100: oled_data = 16'b1011001000101000;
				18'b001010100100011100: oled_data = 16'b1011001000101000;
				18'b001010100110011100: oled_data = 16'b1010101000101000;
				18'b001000011000011101: oled_data = 16'b1010110010100111;
				18'b001000011010011101: oled_data = 16'b1010110010100111;
				18'b001000011100011101: oled_data = 16'b1010110010100111;
				18'b001000011110011101: oled_data = 16'b1010110010101000;
				18'b001000100000011101: oled_data = 16'b1010110010100111;
				18'b001000100010011101: oled_data = 16'b1100010101101011;
				18'b001000100100011101: oled_data = 16'b1101010011010011;
				18'b001000100110011101: oled_data = 16'b1101110010110101;
				18'b001000101000011101: oled_data = 16'b1101110011010110;
				18'b001000101010011101: oled_data = 16'b1101110010110101;
				18'b001000101100011101: oled_data = 16'b1101010010010101;
				18'b001000101110011101: oled_data = 16'b1101110011010110;
				18'b001000110000011101: oled_data = 16'b1101110011010101;
				18'b001000110010011101: oled_data = 16'b1101010001110100;
				18'b001000110100011101: oled_data = 16'b1101110011010110;
				18'b001000110110011101: oled_data = 16'b1101110011010101;
				18'b001000111000011101: oled_data = 16'b1101110011010101;
				18'b001000111010011101: oled_data = 16'b1101110011010101;
				18'b001000111100011101: oled_data = 16'b1101110010110101;
				18'b001000111110011101: oled_data = 16'b1101010001110100;
				18'b001001000000011101: oled_data = 16'b1101110010110101;
				18'b001001000010011101: oled_data = 16'b1101110011010110;
				18'b001001000100011101: oled_data = 16'b1101110011010101;
				18'b001001000110011101: oled_data = 16'b1101010010110101;
				18'b001001001000011101: oled_data = 16'b1110011000111001;
				18'b001001001010011101: oled_data = 16'b1110111100011010;
				18'b001001001100011101: oled_data = 16'b1101111001111000;
				18'b001001001110011101: oled_data = 16'b1101110011010101;
				18'b001001010000011101: oled_data = 16'b1101110011010101;
				18'b001001010010011101: oled_data = 16'b1101110111111000;
				18'b001001010100011101: oled_data = 16'b1101111010011010;
				18'b001001010110011101: oled_data = 16'b1101010011010101;
				18'b001001011000011101: oled_data = 16'b1101010001110100;
				18'b001001011010011101: oled_data = 16'b1101110010110101;
				18'b001001011100011101: oled_data = 16'b1101110011010101;
				18'b001001011110011101: oled_data = 16'b1101110011010101;
				18'b001001100000011101: oled_data = 16'b1101110011010101;
				18'b001001100010011101: oled_data = 16'b1101110011010110;
				18'b001001100100011101: oled_data = 16'b1101010010010100;
				18'b001001100110011101: oled_data = 16'b1101010010010100;
				18'b001001101000011101: oled_data = 16'b1101110100110110;
				18'b001001101010011101: oled_data = 16'b1110011000111001;
				18'b001001101100011101: oled_data = 16'b1101110100010110;
				18'b001001101110011101: oled_data = 16'b0101100111101000;
				18'b001001110000011101: oled_data = 16'b0111101111101111;
				18'b001001110010011101: oled_data = 16'b1110111101111011;
				18'b001001110100011101: oled_data = 16'b1101011001011000;
				18'b001001110110011101: oled_data = 16'b1100110100110101;
				18'b001001111000011101: oled_data = 16'b1110111011111011;
				18'b001001111010011101: oled_data = 16'b1110111100111011;
				18'b001001111100011101: oled_data = 16'b1101111000111001;
				18'b001001111110011101: oled_data = 16'b1010101101101111;
				18'b001010000000011101: oled_data = 16'b1110010011010011;
				18'b001010000010011101: oled_data = 16'b1110010011010011;
				18'b001010000100011101: oled_data = 16'b1011101010001010;
				18'b001010000110011101: oled_data = 16'b1011001000101001;
				18'b001010001000011101: oled_data = 16'b1100001011101011;
				18'b001010001010011101: oled_data = 16'b1100001100101100;
				18'b001010001100011101: oled_data = 16'b1011001000101001;
				18'b001010001110011101: oled_data = 16'b1011101001001001;
				18'b001010010000011101: oled_data = 16'b1011001000101000;
				18'b001010010010011101: oled_data = 16'b1011001001001001;
				18'b001010010100011101: oled_data = 16'b1011101001001001;
				18'b001010010110011101: oled_data = 16'b1010001000001000;
				18'b001010011000011101: oled_data = 16'b1001000101100110;
				18'b001010011010011101: oled_data = 16'b1010101000001000;
				18'b001010011100011101: oled_data = 16'b1011001000101001;
				18'b001010011110011101: oled_data = 16'b1011001000101000;
				18'b001010100000011101: oled_data = 16'b1011001000101001;
				18'b001010100010011101: oled_data = 16'b1011001000101000;
				18'b001010100100011101: oled_data = 16'b1011001000101000;
				18'b001010100110011101: oled_data = 16'b1010101000101000;
				18'b001000011000011110: oled_data = 16'b1010110010100111;
				18'b001000011010011110: oled_data = 16'b1010110010100111;
				18'b001000011100011110: oled_data = 16'b1010110010100111;
				18'b001000011110011110: oled_data = 16'b1010110010100111;
				18'b001000100000011110: oled_data = 16'b1011010011001000;
				18'b001000100010011110: oled_data = 16'b1100110110001101;
				18'b001000100100011110: oled_data = 16'b1100110010010100;
				18'b001000100110011110: oled_data = 16'b1101110011010101;
				18'b001000101000011110: oled_data = 16'b1101110011010110;
				18'b001000101010011110: oled_data = 16'b1101010010010100;
				18'b001000101100011110: oled_data = 16'b1101110011010110;
				18'b001000101110011110: oled_data = 16'b1101110011010101;
				18'b001000110000011110: oled_data = 16'b1101110011010110;
				18'b001000110010011110: oled_data = 16'b1101010001110100;
				18'b001000110100011110: oled_data = 16'b1101110010110101;
				18'b001000110110011110: oled_data = 16'b1101110011010101;
				18'b001000111000011110: oled_data = 16'b1101110011010101;
				18'b001000111010011110: oled_data = 16'b1101110011010110;
				18'b001000111100011110: oled_data = 16'b1101010010010101;
				18'b001000111110011110: oled_data = 16'b1101010001110100;
				18'b001001000000011110: oled_data = 16'b1101110010110101;
				18'b001001000010011110: oled_data = 16'b1101110011010101;
				18'b001001000100011110: oled_data = 16'b1101110010110101;
				18'b001001000110011110: oled_data = 16'b1101010100110110;
				18'b001001001000011110: oled_data = 16'b1110011011011011;
				18'b001001001010011110: oled_data = 16'b1110011100011010;
				18'b001001001100011110: oled_data = 16'b1110011010011001;
				18'b001001001110011110: oled_data = 16'b1101110011110101;
				18'b001001010000011110: oled_data = 16'b1101010011010101;
				18'b001001010010011110: oled_data = 16'b1110011010011010;
				18'b001001010100011110: oled_data = 16'b1101111001011001;
				18'b001001010110011110: oled_data = 16'b1100010001010011;
				18'b001001011000011110: oled_data = 16'b1101010010110101;
				18'b001001011010011110: oled_data = 16'b1101110011010101;
				18'b001001011100011110: oled_data = 16'b1101110011010101;
				18'b001001011110011110: oled_data = 16'b1101110011010101;
				18'b001001100000011110: oled_data = 16'b1101110011010101;
				18'b001001100010011110: oled_data = 16'b1101110011010110;
				18'b001001100100011110: oled_data = 16'b1101010001110100;
				18'b001001100110011110: oled_data = 16'b1101110010110101;
				18'b001001101000011110: oled_data = 16'b1101110110111000;
				18'b001001101010011110: oled_data = 16'b1101010110110111;
				18'b001001101100011110: oled_data = 16'b1100110100010101;
				18'b001001101110011110: oled_data = 16'b0100101000001000;
				18'b001001110000011110: oled_data = 16'b1100011000011000;
				18'b001001110010011110: oled_data = 16'b1110011100111011;
				18'b001001110100011110: oled_data = 16'b1100010111110110;
				18'b001001110110011110: oled_data = 16'b1101011001011000;
				18'b001001111000011110: oled_data = 16'b1101111001111001;
				18'b001001111010011110: oled_data = 16'b1101111010011001;
				18'b001001111100011110: oled_data = 16'b1101111010011010;
				18'b001001111110011110: oled_data = 16'b1100010010010011;
				18'b001010000000011110: oled_data = 16'b1110110100010100;
				18'b001010000010011110: oled_data = 16'b1101001111110000;
				18'b001010000100011110: oled_data = 16'b1011001000101001;
				18'b001010000110011110: oled_data = 16'b1011101001001001;
				18'b001010001000011110: oled_data = 16'b1100001100001100;
				18'b001010001010011110: oled_data = 16'b1011101010001010;
				18'b001010001100011110: oled_data = 16'b1011001001001001;
				18'b001010001110011110: oled_data = 16'b1011001001001001;
				18'b001010010000011110: oled_data = 16'b1010101000101000;
				18'b001010010010011110: oled_data = 16'b1011001001001001;
				18'b001010010100011110: oled_data = 16'b1010101000101000;
				18'b001010010110011110: oled_data = 16'b1000100101100110;
				18'b001010011000011110: oled_data = 16'b1001100110100111;
				18'b001010011010011110: oled_data = 16'b1011101010001010;
				18'b001010011100011110: oled_data = 16'b1011101010101010;
				18'b001010011110011110: oled_data = 16'b1011001000101000;
				18'b001010100000011110: oled_data = 16'b1011001000101001;
				18'b001010100010011110: oled_data = 16'b1011001000101000;
				18'b001010100100011110: oled_data = 16'b1011001000101000;
				18'b001010100110011110: oled_data = 16'b1010101000101000;
				18'b001000011000011111: oled_data = 16'b1011110101001001;
				18'b001000011010011111: oled_data = 16'b1011010100001000;
				18'b001000011100011111: oled_data = 16'b1010110011001000;
				18'b001000011110011111: oled_data = 16'b1010110011101000;
				18'b001000100000011111: oled_data = 16'b1100010110101010;
				18'b001000100010011111: oled_data = 16'b1101010101110000;
				18'b001000100100011111: oled_data = 16'b1101010001110100;
				18'b001000100110011111: oled_data = 16'b1101110010110101;
				18'b001000101000011111: oled_data = 16'b1101010010010101;
				18'b001000101010011111: oled_data = 16'b1101010001110100;
				18'b001000101100011111: oled_data = 16'b1110010011110110;
				18'b001000101110011111: oled_data = 16'b1101110011010110;
				18'b001000110000011111: oled_data = 16'b1101110011010110;
				18'b001000110010011111: oled_data = 16'b1101010010010101;
				18'b001000110100011111: oled_data = 16'b1101110010110101;
				18'b001000110110011111: oled_data = 16'b1101110011010110;
				18'b001000111000011111: oled_data = 16'b1101110011010101;
				18'b001000111010011111: oled_data = 16'b1101110011010101;
				18'b001000111100011111: oled_data = 16'b1101010001110100;
				18'b001000111110011111: oled_data = 16'b1100110001010011;
				18'b001001000000011111: oled_data = 16'b1101110010110101;
				18'b001001000010011111: oled_data = 16'b1101110011010101;
				18'b001001000100011111: oled_data = 16'b1101110010110101;
				18'b001001000110011111: oled_data = 16'b1101110111011000;
				18'b001001001000011111: oled_data = 16'b1110111100011011;
				18'b001001001010011111: oled_data = 16'b1110011100011010;
				18'b001001001100011111: oled_data = 16'b1110011010111001;
				18'b001001001110011111: oled_data = 16'b1101110011110101;
				18'b001001010000011111: oled_data = 16'b1101010100010110;
				18'b001001010010011111: oled_data = 16'b1101111010011001;
				18'b001001010100011111: oled_data = 16'b1101010111110111;
				18'b001001010110011111: oled_data = 16'b1101010011010101;
				18'b001001011000011111: oled_data = 16'b1101110011010110;
				18'b001001011010011111: oled_data = 16'b1101110011010101;
				18'b001001011100011111: oled_data = 16'b1101110011010101;
				18'b001001011110011111: oled_data = 16'b1101110011010101;
				18'b001001100000011111: oled_data = 16'b1101110011010101;
				18'b001001100010011111: oled_data = 16'b1101110010110101;
				18'b001001100100011111: oled_data = 16'b1101010001110100;
				18'b001001100110011111: oled_data = 16'b1101010011110101;
				18'b001001101000011111: oled_data = 16'b1110011010011010;
				18'b001001101010011111: oled_data = 16'b1101111001011001;
				18'b001001101100011111: oled_data = 16'b1011110101010101;
				18'b001001101110011111: oled_data = 16'b0011100110000110;
				18'b001001110000011111: oled_data = 16'b0101101010101010;
				18'b001001110010011111: oled_data = 16'b0101001001101000;
				18'b001001110100011111: oled_data = 16'b0100101000100111;
				18'b001001110110011111: oled_data = 16'b0100001000000110;
				18'b001001111000011111: oled_data = 16'b0011100110000101;
				18'b001001111010011111: oled_data = 16'b0100100111100111;
				18'b001001111100011111: oled_data = 16'b0110001001001001;
				18'b001001111110011111: oled_data = 16'b1100110010110010;
				18'b001010000000011111: oled_data = 16'b1110110100010100;
				18'b001010000010011111: oled_data = 16'b1100001100001101;
				18'b001010000100011111: oled_data = 16'b1011001000101001;
				18'b001010000110011111: oled_data = 16'b1011101001001001;
				18'b001010001000011111: oled_data = 16'b1011101010001010;
				18'b001010001010011111: oled_data = 16'b1011001001001001;
				18'b001010001100011111: oled_data = 16'b1011001001001001;
				18'b001010001110011111: oled_data = 16'b1010101000101000;
				18'b001010010000011111: oled_data = 16'b1011001001001001;
				18'b001010010010011111: oled_data = 16'b1011001000101001;
				18'b001010010100011111: oled_data = 16'b1001000110000111;
				18'b001010010110011111: oled_data = 16'b1001000101100110;
				18'b001010011000011111: oled_data = 16'b1011001001001010;
				18'b001010011010011111: oled_data = 16'b1101001111101111;
				18'b001010011100011111: oled_data = 16'b1011101010001010;
				18'b001010011110011111: oled_data = 16'b1011001000101000;
				18'b001010100000011111: oled_data = 16'b1011001000101001;
				18'b001010100010011111: oled_data = 16'b1011001000101000;
				18'b001010100100011111: oled_data = 16'b1011001000101000;
				18'b001010100110011111: oled_data = 16'b1010101000101000;
				18'b001000011000100000: oled_data = 16'b1101110110001111;
				18'b001000011010100000: oled_data = 16'b1101010110101110;
				18'b001000011100100000: oled_data = 16'b1100110111001100;
				18'b001000011110100000: oled_data = 16'b1100110111001100;
				18'b001000100000100000: oled_data = 16'b1101010111101101;
				18'b001000100010100000: oled_data = 16'b1101010100010010;
				18'b001000100100100000: oled_data = 16'b1101010010010101;
				18'b001000100110100000: oled_data = 16'b1101010010010100;
				18'b001000101000100000: oled_data = 16'b1101110010010101;
				18'b001000101010100000: oled_data = 16'b1101110010110101;
				18'b001000101100100000: oled_data = 16'b1110010011110110;
				18'b001000101110100000: oled_data = 16'b1101110011010110;
				18'b001000110000100000: oled_data = 16'b1101110011010101;
				18'b001000110010100000: oled_data = 16'b1101110010110101;
				18'b001000110100100000: oled_data = 16'b1101010001110100;
				18'b001000110110100000: oled_data = 16'b1101110011010110;
				18'b001000111000100000: oled_data = 16'b1101110011010101;
				18'b001000111010100000: oled_data = 16'b1101110011010101;
				18'b001000111100100000: oled_data = 16'b1101010001010011;
				18'b001000111110100000: oled_data = 16'b1101010011010101;
				18'b001001000000100000: oled_data = 16'b1101110011010101;
				18'b001001000010100000: oled_data = 16'b1101110011010101;
				18'b001001000100100000: oled_data = 16'b1101010011110101;
				18'b001001000110100000: oled_data = 16'b1110111010111010;
				18'b001001001000100000: oled_data = 16'b1110111100011010;
				18'b001001001010100000: oled_data = 16'b1101111011011001;
				18'b001001001100100000: oled_data = 16'b1101011001011000;
				18'b001001001110100000: oled_data = 16'b1100110010010100;
				18'b001001010000100000: oled_data = 16'b1100110011110101;
				18'b001001010010100000: oled_data = 16'b1110011011011010;
				18'b001001010100100000: oled_data = 16'b1110011010011010;
				18'b001001010110100000: oled_data = 16'b1101110011110110;
				18'b001001011000100000: oled_data = 16'b1101110011010110;
				18'b001001011010100000: oled_data = 16'b1101110011010101;
				18'b001001011100100000: oled_data = 16'b1101110011010101;
				18'b001001011110100000: oled_data = 16'b1101110011010101;
				18'b001001100000100000: oled_data = 16'b1101110011010110;
				18'b001001100010100000: oled_data = 16'b1101010001110100;
				18'b001001100100100000: oled_data = 16'b1101010010010101;
				18'b001001100110100000: oled_data = 16'b1101110110110111;
				18'b001001101000100000: oled_data = 16'b1110111100111010;
				18'b001001101010100000: oled_data = 16'b1110111100111011;
				18'b001001101100100000: oled_data = 16'b1100110111110110;
				18'b001001101110100000: oled_data = 16'b0101101010001001;
				18'b001001110000100000: oled_data = 16'b0101001001001001;
				18'b001001110010100000: oled_data = 16'b0101001001101001;
				18'b001001110100100000: oled_data = 16'b0101101010001001;
				18'b001001110110100000: oled_data = 16'b0110001011001010;
				18'b001001111000100000: oled_data = 16'b0111001101001100;
				18'b001001111010100000: oled_data = 16'b0111101110001101;
				18'b001001111100100000: oled_data = 16'b1001110000010000;
				18'b001001111110100000: oled_data = 16'b1101110011010011;
				18'b001010000000100000: oled_data = 16'b1110010011010011;
				18'b001010000010100000: oled_data = 16'b1011001001101010;
				18'b001010000100100000: oled_data = 16'b1011001000101001;
				18'b001010000110100000: oled_data = 16'b1011001001001001;
				18'b001010001000100000: oled_data = 16'b1011001001001001;
				18'b001010001010100000: oled_data = 16'b1011001001001001;
				18'b001010001100100000: oled_data = 16'b1011001001001001;
				18'b001010001110100000: oled_data = 16'b1010101000101001;
				18'b001010010000100000: oled_data = 16'b1011001001001001;
				18'b001010010010100000: oled_data = 16'b1001100110100111;
				18'b001010010100100000: oled_data = 16'b1000100101000110;
				18'b001010010110100000: oled_data = 16'b1010000110101000;
				18'b001010011000100000: oled_data = 16'b1100101101001101;
				18'b001010011010100000: oled_data = 16'b1100001100001100;
				18'b001010011100100000: oled_data = 16'b1011001000101000;
				18'b001010011110100000: oled_data = 16'b1011001000101001;
				18'b001010100000100000: oled_data = 16'b1011001000101001;
				18'b001010100010100000: oled_data = 16'b1011001000101000;
				18'b001010100100100000: oled_data = 16'b1011001000101000;
				18'b001010100110100000: oled_data = 16'b1010101000101000;
				18'b001000011000100001: oled_data = 16'b1101110011010110;
				18'b001000011010100001: oled_data = 16'b1101110011010110;
				18'b001000011100100001: oled_data = 16'b1101110011010101;
				18'b001000011110100001: oled_data = 16'b1101110011010100;
				18'b001000100000100001: oled_data = 16'b1101110011010101;
				18'b001000100010100001: oled_data = 16'b1101010010010101;
				18'b001000100100100001: oled_data = 16'b1101010010010101;
				18'b001000100110100001: oled_data = 16'b1101010010010101;
				18'b001000101000100001: oled_data = 16'b1101110010010101;
				18'b001000101010100001: oled_data = 16'b1101110011010101;
				18'b001000101100100001: oled_data = 16'b1110010011110110;
				18'b001000101110100001: oled_data = 16'b1101110011010110;
				18'b001000110000100001: oled_data = 16'b1101110011010110;
				18'b001000110010100001: oled_data = 16'b1101110011010110;
				18'b001000110100100001: oled_data = 16'b1101110010110101;
				18'b001000110110100001: oled_data = 16'b1101110011010110;
				18'b001000111000100001: oled_data = 16'b1101110011010110;
				18'b001000111010100001: oled_data = 16'b1101110010110101;
				18'b001000111100100001: oled_data = 16'b1101010010010100;
				18'b001000111110100001: oled_data = 16'b1110010101110111;
				18'b001001000000100001: oled_data = 16'b1101110011010110;
				18'b001001000010100001: oled_data = 16'b1101110010110101;
				18'b001001000100100001: oled_data = 16'b1101010110010110;
				18'b001001000110100001: oled_data = 16'b1110111100011011;
				18'b001001001000100001: oled_data = 16'b1110111011111010;
				18'b001001001010100001: oled_data = 16'b1110111011111010;
				18'b001001001100100001: oled_data = 16'b1110011011111010;
				18'b001001001110100001: oled_data = 16'b1101010100110101;
				18'b001001010000100001: oled_data = 16'b1101110110010111;
				18'b001001010010100001: oled_data = 16'b1111011100111011;
				18'b001001010100100001: oled_data = 16'b1110011010011010;
				18'b001001010110100001: oled_data = 16'b1101010011110110;
				18'b001001011000100001: oled_data = 16'b1101110011010110;
				18'b001001011010100001: oled_data = 16'b1101110011010101;
				18'b001001011100100001: oled_data = 16'b1101110011010101;
				18'b001001011110100001: oled_data = 16'b1101110011010101;
				18'b001001100000100001: oled_data = 16'b1101110010110101;
				18'b001001100010100001: oled_data = 16'b1101010001110100;
				18'b001001100100100001: oled_data = 16'b1101010100010101;
				18'b001001100110100001: oled_data = 16'b1110011011011010;
				18'b001001101000100001: oled_data = 16'b1110111100011010;
				18'b001001101010100001: oled_data = 16'b1110011100011010;
				18'b001001101100100001: oled_data = 16'b1110111100011011;
				18'b001001101110100001: oled_data = 16'b1110011011111010;
				18'b001001110000100001: oled_data = 16'b1110011011111010;
				18'b001001110010100001: oled_data = 16'b1110011011111010;
				18'b001001110100100001: oled_data = 16'b1110011011111010;
				18'b001001110110100001: oled_data = 16'b1110111100011010;
				18'b001001111000100001: oled_data = 16'b1110111100011011;
				18'b001001111010100001: oled_data = 16'b1101111011011010;
				18'b001001111100100001: oled_data = 16'b1110011000111000;
				18'b001001111110100001: oled_data = 16'b1110010100010100;
				18'b001010000000100001: oled_data = 16'b1101110001110001;
				18'b001010000010100001: oled_data = 16'b1011001000101001;
				18'b001010000100100001: oled_data = 16'b1011001001001001;
				18'b001010000110100001: oled_data = 16'b1011001001001001;
				18'b001010001000100001: oled_data = 16'b1011001001001001;
				18'b001010001010100001: oled_data = 16'b1011001001001001;
				18'b001010001100100001: oled_data = 16'b1010101000101001;
				18'b001010001110100001: oled_data = 16'b1011001001001001;
				18'b001010010000100001: oled_data = 16'b1010100111101000;
				18'b001010010010100001: oled_data = 16'b1000100101000110;
				18'b001010010100100001: oled_data = 16'b1001000110000111;
				18'b001010010110100001: oled_data = 16'b1011001001101010;
				18'b001010011000100001: oled_data = 16'b1011001010001010;
				18'b001010011010100001: oled_data = 16'b1011001000101001;
				18'b001010011100100001: oled_data = 16'b1011001000101001;
				18'b001010011110100001: oled_data = 16'b1011001000101001;
				18'b001010100000100001: oled_data = 16'b1011001000101001;
				18'b001010100010100001: oled_data = 16'b1011001000101000;
				18'b001010100100100001: oled_data = 16'b1011001000101000;
				18'b001010100110100001: oled_data = 16'b1010101000101000;
				18'b001000011000100010: oled_data = 16'b1101110011010110;
				18'b001000011010100010: oled_data = 16'b1101110011010110;
				18'b001000011100100010: oled_data = 16'b1101110011010110;
				18'b001000011110100010: oled_data = 16'b1101110011010110;
				18'b001000100000100010: oled_data = 16'b1101110011010110;
				18'b001000100010100010: oled_data = 16'b1101010010010101;
				18'b001000100100100010: oled_data = 16'b1100110001010100;
				18'b001000100110100010: oled_data = 16'b1101110010110101;
				18'b001000101000100010: oled_data = 16'b1101010001110100;
				18'b001000101010100010: oled_data = 16'b1101110011010110;
				18'b001000101100100010: oled_data = 16'b1101010010010100;
				18'b001000101110100010: oled_data = 16'b1101110011010101;
				18'b001000110000100010: oled_data = 16'b1101110011010101;
				18'b001000110010100010: oled_data = 16'b1101110011010101;
				18'b001000110100100010: oled_data = 16'b1101110011010110;
				18'b001000110110100010: oled_data = 16'b1101110011010101;
				18'b001000111000100010: oled_data = 16'b1110010011010110;
				18'b001000111010100010: oled_data = 16'b1101110010010101;
				18'b001000111100100010: oled_data = 16'b1101010011110101;
				18'b001000111110100010: oled_data = 16'b1101111000011001;
				18'b001001000000100010: oled_data = 16'b1101110011010101;
				18'b001001000010100010: oled_data = 16'b1101010011010101;
				18'b001001000100100010: oled_data = 16'b1110011010011010;
				18'b001001000110100010: oled_data = 16'b1110111100011010;
				18'b001001001000100010: oled_data = 16'b1110111011111010;
				18'b001001001010100010: oled_data = 16'b1110111011111010;
				18'b001001001100100010: oled_data = 16'b1110111100011010;
				18'b001001001110100010: oled_data = 16'b1100110110010101;
				18'b001001010000100010: oled_data = 16'b1101111000111000;
				18'b001001010010100010: oled_data = 16'b1110111100111011;
				18'b001001010100100010: oled_data = 16'b1110011010111010;
				18'b001001010110100010: oled_data = 16'b1101010011110110;
				18'b001001011000100010: oled_data = 16'b1101110011010110;
				18'b001001011010100010: oled_data = 16'b1101110011010101;
				18'b001001011100100010: oled_data = 16'b1101110011010101;
				18'b001001011110100010: oled_data = 16'b1101110011010110;
				18'b001001100000100010: oled_data = 16'b1101010010010100;
				18'b001001100010100010: oled_data = 16'b1101010010110100;
				18'b001001100100100010: oled_data = 16'b1110011001011000;
				18'b001001100110100010: oled_data = 16'b1110011100111011;
				18'b001001101000100010: oled_data = 16'b1110111100011010;
				18'b001001101010100010: oled_data = 16'b1110111100011010;
				18'b001001101100100010: oled_data = 16'b1110111100011010;
				18'b001001101110100010: oled_data = 16'b1110111100011010;
				18'b001001110000100010: oled_data = 16'b1110111100011010;
				18'b001001110010100010: oled_data = 16'b1110111100011010;
				18'b001001110100100010: oled_data = 16'b1110111100011010;
				18'b001001110110100010: oled_data = 16'b1110111100011010;
				18'b001001111000100010: oled_data = 16'b1101111010111001;
				18'b001001111010100010: oled_data = 16'b1110011011111001;
				18'b001001111100100010: oled_data = 16'b1101110110110110;
				18'b001001111110100010: oled_data = 16'b1110110100010100;
				18'b001010000000100010: oled_data = 16'b1100101111001111;
				18'b001010000010100010: oled_data = 16'b1010101000001000;
				18'b001010000100100010: oled_data = 16'b1011101001001001;
				18'b001010000110100010: oled_data = 16'b1011001001001001;
				18'b001010001000100010: oled_data = 16'b1011001001001001;
				18'b001010001010100010: oled_data = 16'b1011001001001001;
				18'b001010001100100010: oled_data = 16'b1010101000101000;
				18'b001010001110100010: oled_data = 16'b1011001001001001;
				18'b001010010000100010: oled_data = 16'b1001000101100110;
				18'b001010010010100010: oled_data = 16'b1000100101100110;
				18'b001010010100100010: oled_data = 16'b1010100111101000;
				18'b001010010110100010: oled_data = 16'b1011110011010011;
				18'b001010011000100010: oled_data = 16'b1011001100001100;
				18'b001010011010100010: oled_data = 16'b1011001000101000;
				18'b001010011100100010: oled_data = 16'b1011001001001001;
				18'b001010011110100010: oled_data = 16'b1011001001001001;
				18'b001010100000100010: oled_data = 16'b1011001000101001;
				18'b001010100010100010: oled_data = 16'b1011001000101000;
				18'b001010100100100010: oled_data = 16'b1010101000101000;
				18'b001010100110100010: oled_data = 16'b1010101000101000;
				18'b001000011000100011: oled_data = 16'b1101110011010110;
				18'b001000011010100011: oled_data = 16'b1101110011010110;
				18'b001000011100100011: oled_data = 16'b1101110011010110;
				18'b001000011110100011: oled_data = 16'b1101110011010110;
				18'b001000100000100011: oled_data = 16'b1101110011010110;
				18'b001000100010100011: oled_data = 16'b1101010001110100;
				18'b001000100100100011: oled_data = 16'b1100110000110011;
				18'b001000100110100011: oled_data = 16'b1101110010110101;
				18'b001000101000100011: oled_data = 16'b1101010001110100;
				18'b001000101010100011: oled_data = 16'b1101110011010101;
				18'b001000101100100011: oled_data = 16'b1101010001110100;
				18'b001000101110100011: oled_data = 16'b1101110011010110;
				18'b001000110000100011: oled_data = 16'b1101110011010101;
				18'b001000110010100011: oled_data = 16'b1110010011010101;
				18'b001000110100100011: oled_data = 16'b1110010011010101;
				18'b001000110110100011: oled_data = 16'b1110010011010101;
				18'b001000111000100011: oled_data = 16'b1110010011010101;
				18'b001000111010100011: oled_data = 16'b1101010001110100;
				18'b001000111100100011: oled_data = 16'b1101010100110110;
				18'b001000111110100011: oled_data = 16'b1110011001011001;
				18'b001001000000100011: oled_data = 16'b1101110010110101;
				18'b001001000010100011: oled_data = 16'b1101110101110111;
				18'b001001000100100011: oled_data = 16'b1110111100011011;
				18'b001001000110100011: oled_data = 16'b1110011100011010;
				18'b001001001000100011: oled_data = 16'b1110111100111011;
				18'b001001001010100011: oled_data = 16'b1110111100111011;
				18'b001001001100100011: oled_data = 16'b1110111101011011;
				18'b001001001110100011: oled_data = 16'b1101011000010111;
				18'b001001010000100011: oled_data = 16'b1110011010111010;
				18'b001001010010100011: oled_data = 16'b1110111101011011;
				18'b001001010100100011: oled_data = 16'b1110011011011010;
				18'b001001010110100011: oled_data = 16'b1101010100010110;
				18'b001001011000100011: oled_data = 16'b1110010011110110;
				18'b001001011010100011: oled_data = 16'b1110010011110110;
				18'b001001011100100011: oled_data = 16'b1101110011110110;
				18'b001001011110100011: oled_data = 16'b1101110011010101;
				18'b001001100000100011: oled_data = 16'b1101010001010100;
				18'b001001100010100011: oled_data = 16'b1101110101010110;
				18'b001001100100100011: oled_data = 16'b1110111100011011;
				18'b001001100110100011: oled_data = 16'b1110011100011011;
				18'b001001101000100011: oled_data = 16'b1110111100011010;
				18'b001001101010100011: oled_data = 16'b1110111100011010;
				18'b001001101100100011: oled_data = 16'b1110111100011010;
				18'b001001101110100011: oled_data = 16'b1110111100011010;
				18'b001001110000100011: oled_data = 16'b1110111100011010;
				18'b001001110010100011: oled_data = 16'b1110011100011010;
				18'b001001110100100011: oled_data = 16'b1110111100011010;
				18'b001001110110100011: oled_data = 16'b1110011011111010;
				18'b001001111000100011: oled_data = 16'b1101111010011000;
				18'b001001111010100011: oled_data = 16'b1110111100111010;
				18'b001001111100100011: oled_data = 16'b1101010110010101;
				18'b001001111110100011: oled_data = 16'b1110110100010100;
				18'b001010000000100011: oled_data = 16'b1100001100101100;
				18'b001010000010100011: oled_data = 16'b1010101000101001;
				18'b001010000100100011: oled_data = 16'b1011101001001001;
				18'b001010000110100011: oled_data = 16'b1011001001001001;
				18'b001010001000100011: oled_data = 16'b1011001001001001;
				18'b001010001010100011: oled_data = 16'b1011001000101001;
				18'b001010001100100011: oled_data = 16'b1010101000101001;
				18'b001010001110100011: oled_data = 16'b1010000111101000;
				18'b001010010000100011: oled_data = 16'b1000100101000110;
				18'b001010010010100011: oled_data = 16'b1001100111000111;
				18'b001010010100100011: oled_data = 16'b1011001011101100;
				18'b001010010110100011: oled_data = 16'b1100011010111010;
				18'b001010011000100011: oled_data = 16'b1011010010110011;
				18'b001010011010100011: oled_data = 16'b1011001000001000;
				18'b001010011100100011: oled_data = 16'b1011001000101001;
				18'b001010011110100011: oled_data = 16'b1011001000101001;
				18'b001010100000100011: oled_data = 16'b1011001000101001;
				18'b001010100010100011: oled_data = 16'b1011001000101000;
				18'b001010100100100011: oled_data = 16'b1010101000101000;
				18'b001010100110100011: oled_data = 16'b1010101000101000;
				18'b001000011000100100: oled_data = 16'b1101110011010101;
				18'b001000011010100100: oled_data = 16'b1101110011010110;
				18'b001000011100100100: oled_data = 16'b1101110011010101;
				18'b001000011110100100: oled_data = 16'b1101110011010110;
				18'b001000100000100100: oled_data = 16'b1101110011010110;
				18'b001000100010100100: oled_data = 16'b1100110000110011;
				18'b001000100100100100: oled_data = 16'b1100110001010100;
				18'b001000100110100100: oled_data = 16'b1101010010010101;
				18'b001000101000100100: oled_data = 16'b1101010010010101;
				18'b001000101010100100: oled_data = 16'b1101110010110101;
				18'b001000101100100100: oled_data = 16'b1101010010010101;
				18'b001000101110100100: oled_data = 16'b1101110011010110;
				18'b001000110000100100: oled_data = 16'b1101110011010110;
				18'b001000110010100100: oled_data = 16'b1101110011010110;
				18'b001000110100100100: oled_data = 16'b1101110011010110;
				18'b001000110110100100: oled_data = 16'b1101110011010110;
				18'b001000111000100100: oled_data = 16'b1101110011010110;
				18'b001000111010100100: oled_data = 16'b1101010001110100;
				18'b001000111100100100: oled_data = 16'b1101110110010111;
				18'b001000111110100100: oled_data = 16'b1110011001111001;
				18'b001001000000100100: oled_data = 16'b1101010011010100;
				18'b001001000010100100: oled_data = 16'b1110011010011001;
				18'b001001000100100100: oled_data = 16'b1110111100011010;
				18'b001001000110100100: oled_data = 16'b1110011011011001;
				18'b001001001000100100: oled_data = 16'b1010110101010011;
				18'b001001001010100100: oled_data = 16'b1001110011010010;
				18'b001001001100100100: oled_data = 16'b1011010101110101;
				18'b001001001110100100: oled_data = 16'b1011010101110101;
				18'b001001010000100100: oled_data = 16'b1100010111010110;
				18'b001001010010100100: oled_data = 16'b1100111000110111;
				18'b001001010100100100: oled_data = 16'b1100010111110110;
				18'b001001010110100100: oled_data = 16'b1011110010010100;
				18'b001001011000100100: oled_data = 16'b1100110010110100;
				18'b001001011010100100: oled_data = 16'b1100110010110100;
				18'b001001011100100100: oled_data = 16'b1101010011010101;
				18'b001001011110100100: oled_data = 16'b1100110010010100;
				18'b001001100000100100: oled_data = 16'b1101010011110101;
				18'b001001100010100100: oled_data = 16'b1110011010111011;
				18'b001001100100100100: oled_data = 16'b1110111100011011;
				18'b001001100110100100: oled_data = 16'b1110011100011011;
				18'b001001101000100100: oled_data = 16'b1110111100011010;
				18'b001001101010100100: oled_data = 16'b1110111100011010;
				18'b001001101100100100: oled_data = 16'b1110111100011010;
				18'b001001101110100100: oled_data = 16'b1110111100011010;
				18'b001001110000100100: oled_data = 16'b1110111100011010;
				18'b001001110010100100: oled_data = 16'b1110111100011010;
				18'b001001110100100100: oled_data = 16'b1110111100011010;
				18'b001001110110100100: oled_data = 16'b1101111010011000;
				18'b001001111000100100: oled_data = 16'b1110011011111010;
				18'b001001111010100100: oled_data = 16'b1110011100011010;
				18'b001001111100100100: oled_data = 16'b1101010101010100;
				18'b001001111110100100: oled_data = 16'b1110110011110011;
				18'b001010000000100100: oled_data = 16'b1011001010101011;
				18'b001010000010100100: oled_data = 16'b1011001000101001;
				18'b001010000100100100: oled_data = 16'b1011001001001001;
				18'b001010000110100100: oled_data = 16'b1011001001001001;
				18'b001010001000100100: oled_data = 16'b1011001001001001;
				18'b001010001010100100: oled_data = 16'b1010101000101000;
				18'b001010001100100100: oled_data = 16'b1011001000101001;
				18'b001010001110100100: oled_data = 16'b1001000101100110;
				18'b001010010000100100: oled_data = 16'b1001000101100111;
				18'b001010010010100100: oled_data = 16'b1010101000001001;
				18'b001010010100100100: oled_data = 16'b1011110010110011;
				18'b001010010110100100: oled_data = 16'b1011111100111100;
				18'b001010011000100100: oled_data = 16'b1011111001011001;
				18'b001010011010100100: oled_data = 16'b1011001010001010;
				18'b001010011100100100: oled_data = 16'b1011101001001001;
				18'b001010011110100100: oled_data = 16'b1011001001001001;
				18'b001010100000100100: oled_data = 16'b1011001000101001;
				18'b001010100010100100: oled_data = 16'b1011001000101000;
				18'b001010100100100100: oled_data = 16'b1010101000101000;
				18'b001010100110100100: oled_data = 16'b1010101000101000;
				18'b001000011000100101: oled_data = 16'b1101110011010101;
				18'b001000011010100101: oled_data = 16'b1101110011010110;
				18'b001000011100100101: oled_data = 16'b1101110011010110;
				18'b001000011110100101: oled_data = 16'b1101110011010110;
				18'b001000100000100101: oled_data = 16'b1101110011010110;
				18'b001000100010100101: oled_data = 16'b1101010001010100;
				18'b001000100100100101: oled_data = 16'b1101110010110101;
				18'b001000100110100101: oled_data = 16'b1100110000110011;
				18'b001000101000100101: oled_data = 16'b1101010010010101;
				18'b001000101010100101: oled_data = 16'b1101010010010101;
				18'b001000101100100101: oled_data = 16'b1101110010110101;
				18'b001000101110100101: oled_data = 16'b1101110011010110;
				18'b001000110000100101: oled_data = 16'b1101110011010101;
				18'b001000110010100101: oled_data = 16'b1101110011010101;
				18'b001000110100100101: oled_data = 16'b1101110011010101;
				18'b001000110110100101: oled_data = 16'b1101110011010101;
				18'b001000111000100101: oled_data = 16'b1101110011010101;
				18'b001000111010100101: oled_data = 16'b1101010001110100;
				18'b001000111100100101: oled_data = 16'b1101111000011001;
				18'b001000111110100101: oled_data = 16'b1110011001111001;
				18'b001001000000100101: oled_data = 16'b1101010110110110;
				18'b001001000010100101: oled_data = 16'b1110111011111010;
				18'b001001000100100101: oled_data = 16'b1110111100011010;
				18'b001001000110100101: oled_data = 16'b1100111000110111;
				18'b001001001000100101: oled_data = 16'b0100101000000111;
				18'b001001001010100101: oled_data = 16'b0010000011100011;
				18'b001001001100100101: oled_data = 16'b0010100100100100;
				18'b001001001110100101: oled_data = 16'b0011000101000100;
				18'b001001010000100101: oled_data = 16'b0011000101100101;
				18'b001001010010100101: oled_data = 16'b0011100110000101;
				18'b001001010100100101: oled_data = 16'b0011100110000101;
				18'b001001010110100101: oled_data = 16'b0101000111001000;
				18'b001001011000100101: oled_data = 16'b0110001000001001;
				18'b001001011010100101: oled_data = 16'b0110101000001001;
				18'b001001011100100101: oled_data = 16'b0110101001001010;
				18'b001001011110100101: oled_data = 16'b1011110010010011;
				18'b001001100000100101: oled_data = 16'b1110011001111010;
				18'b001001100010100101: oled_data = 16'b1110111100011100;
				18'b001001100100100101: oled_data = 16'b1110011100011011;
				18'b001001100110100101: oled_data = 16'b1110011100011011;
				18'b001001101000100101: oled_data = 16'b1110111100011010;
				18'b001001101010100101: oled_data = 16'b1110111100011010;
				18'b001001101100100101: oled_data = 16'b1110111100011010;
				18'b001001101110100101: oled_data = 16'b1110111100011010;
				18'b001001110000100101: oled_data = 16'b1110111100011010;
				18'b001001110010100101: oled_data = 16'b1110111100011010;
				18'b001001110100100101: oled_data = 16'b1101111010111001;
				18'b001001110110100101: oled_data = 16'b1101111011011001;
				18'b001001111000100101: oled_data = 16'b1110111100011010;
				18'b001001111010100101: oled_data = 16'b1110011010011001;
				18'b001001111100100101: oled_data = 16'b1101010011110011;
				18'b001001111110100101: oled_data = 16'b1110010011010011;
				18'b001010000000100101: oled_data = 16'b1011001001101001;
				18'b001010000010100101: oled_data = 16'b1011001001001001;
				18'b001010000100100101: oled_data = 16'b1011001001001001;
				18'b001010000110100101: oled_data = 16'b1011001001001001;
				18'b001010001000100101: oled_data = 16'b1011101010101010;
				18'b001010001010100101: oled_data = 16'b1011001010001001;
				18'b001010001100100101: oled_data = 16'b1010000111101000;
				18'b001010001110100101: oled_data = 16'b1000100101000110;
				18'b001010010000100101: oled_data = 16'b1010000111101000;
				18'b001010010010100101: oled_data = 16'b1011001010001011;
				18'b001010010100100101: oled_data = 16'b1011111000011000;
				18'b001010010110100101: oled_data = 16'b1011111100011100;
				18'b001010011000100101: oled_data = 16'b1011111100011100;
				18'b001010011010100101: oled_data = 16'b1011110000110000;
				18'b001010011100100101: oled_data = 16'b1011101001101010;
				18'b001010011110100101: oled_data = 16'b1011001001001001;
				18'b001010100000100101: oled_data = 16'b1011001000101001;
				18'b001010100010100101: oled_data = 16'b1011001000101000;
				18'b001010100100100101: oled_data = 16'b1010101000101000;
				18'b001010100110100101: oled_data = 16'b1010101000101000;
				18'b001000011000100110: oled_data = 16'b1101110011010101;
				18'b001000011010100110: oled_data = 16'b1101110011010110;
				18'b001000011100100110: oled_data = 16'b1101110011010110;
				18'b001000011110100110: oled_data = 16'b1101110011010110;
				18'b001000100000100110: oled_data = 16'b1101110011010101;
				18'b001000100010100110: oled_data = 16'b1101010010010100;
				18'b001000100100100110: oled_data = 16'b1101110010110101;
				18'b001000100110100110: oled_data = 16'b1011101111010001;
				18'b001000101000100110: oled_data = 16'b1101110011010101;
				18'b001000101010100110: oled_data = 16'b1100110001010011;
				18'b001000101100100110: oled_data = 16'b1101110010110101;
				18'b001000101110100110: oled_data = 16'b1101110011010101;
				18'b001000110000100110: oled_data = 16'b1101110011010101;
				18'b001000110010100110: oled_data = 16'b1101110011010101;
				18'b001000110100100110: oled_data = 16'b1101110011010101;
				18'b001000110110100110: oled_data = 16'b1101110011010101;
				18'b001000111000100110: oled_data = 16'b1101110011010101;
				18'b001000111010100110: oled_data = 16'b1101010001110100;
				18'b001000111100100110: oled_data = 16'b1110011001111010;
				18'b001000111110100110: oled_data = 16'b1110011011111010;
				18'b001001000000100110: oled_data = 16'b1110011011111010;
				18'b001001000010100110: oled_data = 16'b1110111100011010;
				18'b001001000100100110: oled_data = 16'b1110111100011010;
				18'b001001000110100110: oled_data = 16'b1101011010011001;
				18'b001001001000100110: oled_data = 16'b1010010011110011;
				18'b001001001010100110: oled_data = 16'b1000001111101111;
				18'b001001001100100110: oled_data = 16'b0110101100101100;
				18'b001001001110100110: oled_data = 16'b0101101010101010;
				18'b001001010000100110: oled_data = 16'b0101001001101001;
				18'b001001010010100110: oled_data = 16'b0101001000101000;
				18'b001001010100100110: oled_data = 16'b0100101000101000;
				18'b001001010110100110: oled_data = 16'b0110001001001001;
				18'b001001011000100110: oled_data = 16'b0110001000101001;
				18'b001001011010100110: oled_data = 16'b0101100111101000;
				18'b001001011100100110: oled_data = 16'b0111101011101100;
				18'b001001011110100110: oled_data = 16'b1101111000111001;
				18'b001001100000100110: oled_data = 16'b1110111100111011;
				18'b001001100010100110: oled_data = 16'b1110111100011010;
				18'b001001100100100110: oled_data = 16'b1110011100011011;
				18'b001001100110100110: oled_data = 16'b1110011100011011;
				18'b001001101000100110: oled_data = 16'b1110111100011010;
				18'b001001101010100110: oled_data = 16'b1110111100011010;
				18'b001001101100100110: oled_data = 16'b1110111100011010;
				18'b001001101110100110: oled_data = 16'b1110111100011010;
				18'b001001110000100110: oled_data = 16'b1110111100011010;
				18'b001001110010100110: oled_data = 16'b1110011011111010;
				18'b001001110100100110: oled_data = 16'b1101111010011001;
				18'b001001110110100110: oled_data = 16'b1110111100011010;
				18'b001001111000100110: oled_data = 16'b1110111100111011;
				18'b001001111010100110: oled_data = 16'b1100010100110100;
				18'b001001111100100110: oled_data = 16'b1100110010010011;
				18'b001001111110100110: oled_data = 16'b1101110001110001;
				18'b001010000000100110: oled_data = 16'b1010101000101001;
				18'b001010000010100110: oled_data = 16'b1011001001001001;
				18'b001010000100100110: oled_data = 16'b1011001010101010;
				18'b001010000110100110: oled_data = 16'b1101010000110000;
				18'b001010001000100110: oled_data = 16'b1110010011010011;
				18'b001010001010100110: oled_data = 16'b1100101110101111;
				18'b001010001100100110: oled_data = 16'b1010000111101000;
				18'b001010001110100110: oled_data = 16'b1001100110000111;
				18'b001010010000100110: oled_data = 16'b1011001000001001;
				18'b001010010010100110: oled_data = 16'b1011010000110000;
				18'b001010010100100110: oled_data = 16'b1011111100011100;
				18'b001010010110100110: oled_data = 16'b1011111011111011;
				18'b001010011000100110: oled_data = 16'b1011111100011100;
				18'b001010011010100110: oled_data = 16'b1011110111110111;
				18'b001010011100100110: oled_data = 16'b1011001001001001;
				18'b001010011110100110: oled_data = 16'b1011001000101000;
				18'b001010100000100110: oled_data = 16'b1011001000101001;
				18'b001010100010100110: oled_data = 16'b1011001000101000;
				18'b001010100100100110: oled_data = 16'b1010101000101000;
				18'b001010100110100110: oled_data = 16'b1010101000101000;
				18'b001000011000100111: oled_data = 16'b1101110011010101;
				18'b001000011010100111: oled_data = 16'b1101110011010101;
				18'b001000011100100111: oled_data = 16'b1101110011010110;
				18'b001000011110100111: oled_data = 16'b1101110011010110;
				18'b001000100000100111: oled_data = 16'b1101010010010101;
				18'b001000100010100111: oled_data = 16'b1101010010010100;
				18'b001000100100100111: oled_data = 16'b1100110001010011;
				18'b001000100110100111: oled_data = 16'b1011101111010001;
				18'b001000101000100111: oled_data = 16'b1101110011010101;
				18'b001000101010100111: oled_data = 16'b1100010000010010;
				18'b001000101100100111: oled_data = 16'b1101110011010101;
				18'b001000101110100111: oled_data = 16'b1101110011010101;
				18'b001000110000100111: oled_data = 16'b1101110011010101;
				18'b001000110010100111: oled_data = 16'b1101110011010101;
				18'b001000110100100111: oled_data = 16'b1101110011010101;
				18'b001000110110100111: oled_data = 16'b1101110011010110;
				18'b001000111000100111: oled_data = 16'b1101110010110101;
				18'b001000111010100111: oled_data = 16'b1101010010010100;
				18'b001000111100100111: oled_data = 16'b1110011010111010;
				18'b001000111110100111: oled_data = 16'b1110011100011011;
				18'b001001000000100111: oled_data = 16'b1110111100011010;
				18'b001001000010100111: oled_data = 16'b1110111100011010;
				18'b001001000100100111: oled_data = 16'b1110011100011010;
				18'b001001000110100111: oled_data = 16'b1110111100011011;
				18'b001001001000100111: oled_data = 16'b1110111100111011;
				18'b001001001010100111: oled_data = 16'b1110111100111100;
				18'b001001001100100111: oled_data = 16'b1110111100111011;
				18'b001001001110100111: oled_data = 16'b1110011100011011;
				18'b001001010000100111: oled_data = 16'b1110011011011010;
				18'b001001010010100111: oled_data = 16'b1101111011011010;
				18'b001001010100100111: oled_data = 16'b1110011011111010;
				18'b001001010110100111: oled_data = 16'b1011010011110100;
				18'b001001011000100111: oled_data = 16'b0101101000101001;
				18'b001001011010100111: oled_data = 16'b0101001000001000;
				18'b001001011100100111: oled_data = 16'b1100110110110111;
				18'b001001011110100111: oled_data = 16'b1111011100011100;
				18'b001001100000100111: oled_data = 16'b1110111100011010;
				18'b001001100010100111: oled_data = 16'b1110111100011010;
				18'b001001100100100111: oled_data = 16'b1110011100011010;
				18'b001001100110100111: oled_data = 16'b1110011100011010;
				18'b001001101000100111: oled_data = 16'b1110111100011010;
				18'b001001101010100111: oled_data = 16'b1110111100011010;
				18'b001001101100100111: oled_data = 16'b1110111100011010;
				18'b001001101110100111: oled_data = 16'b1110111100011010;
				18'b001001110000100111: oled_data = 16'b1110111100011010;
				18'b001001110010100111: oled_data = 16'b1101111010011000;
				18'b001001110100100111: oled_data = 16'b1110111100011010;
				18'b001001110110100111: oled_data = 16'b1110111100111011;
				18'b001001111000100111: oled_data = 16'b1101111001011000;
				18'b001001111010100111: oled_data = 16'b1011001111110001;
				18'b001001111100100111: oled_data = 16'b1101110010110100;
				18'b001001111110100111: oled_data = 16'b1101010000110000;
				18'b001010000000100111: oled_data = 16'b1010101000101000;
				18'b001010000010100111: oled_data = 16'b1011001001001001;
				18'b001010000100100111: oled_data = 16'b1101010001010001;
				18'b001010000110100111: oled_data = 16'b1110010011110011;
				18'b001010001000100111: oled_data = 16'b1100001100001101;
				18'b001010001010100111: oled_data = 16'b1011001000101001;
				18'b001010001100100111: oled_data = 16'b1011001000101001;
				18'b001010001110100111: oled_data = 16'b1011001000101001;
				18'b001010010000100111: oled_data = 16'b1011001001101010;
				18'b001010010010100111: oled_data = 16'b1100010111010111;
				18'b001010010100100111: oled_data = 16'b1011111100011100;
				18'b001010010110100111: oled_data = 16'b1011111011111011;
				18'b001010011000100111: oled_data = 16'b1011111011111100;
				18'b001010011010100111: oled_data = 16'b1011111011111100;
				18'b001010011100100111: oled_data = 16'b1011001110001110;
				18'b001010011110100111: oled_data = 16'b1011001000001000;
				18'b001010100000100111: oled_data = 16'b1011001000101001;
				18'b001010100010100111: oled_data = 16'b1010101000101000;
				18'b001010100100100111: oled_data = 16'b1010000111101000;
				18'b001010100110100111: oled_data = 16'b1010101000001000;
				18'b001000011000101000: oled_data = 16'b1101110011010101;
				18'b001000011010101000: oled_data = 16'b1101110011010101;
				18'b001000011100101000: oled_data = 16'b1101110011010101;
				18'b001000011110101000: oled_data = 16'b1101110011010101;
				18'b001000100000101000: oled_data = 16'b1101010001110100;
				18'b001000100010101000: oled_data = 16'b1101010001110100;
				18'b001000100100101000: oled_data = 16'b1011101110110001;
				18'b001000100110101000: oled_data = 16'b1100010000110010;
				18'b001000101000101000: oled_data = 16'b1101110011010101;
				18'b001000101010101000: oled_data = 16'b1100010000110011;
				18'b001000101100101000: oled_data = 16'b1101110011110110;
				18'b001000101110101000: oled_data = 16'b1101110011010101;
				18'b001000110000101000: oled_data = 16'b1101110011010101;
				18'b001000110010101000: oled_data = 16'b1101110011010101;
				18'b001000110100101000: oled_data = 16'b1101110011010101;
				18'b001000110110101000: oled_data = 16'b1101110011010110;
				18'b001000111000101000: oled_data = 16'b1101110010110101;
				18'b001000111010101000: oled_data = 16'b1100110011010101;
				18'b001000111100101000: oled_data = 16'b1110011011011010;
				18'b001000111110101000: oled_data = 16'b1110011100011010;
				18'b001001000000101000: oled_data = 16'b1110111100011010;
				18'b001001000010101000: oled_data = 16'b1110111100011010;
				18'b001001000100101000: oled_data = 16'b1110111100011010;
				18'b001001000110101000: oled_data = 16'b1110111100011010;
				18'b001001001000101000: oled_data = 16'b1110111100011010;
				18'b001001001010101000: oled_data = 16'b1110111100011010;
				18'b001001001100101000: oled_data = 16'b1110111100011010;
				18'b001001001110101000: oled_data = 16'b1110111100011010;
				18'b001001010000101000: oled_data = 16'b1110111100011010;
				18'b001001010010101000: oled_data = 16'b1110111100111011;
				18'b001001010100101000: oled_data = 16'b1101111010111010;
				18'b001001010110101000: oled_data = 16'b0110101010101010;
				18'b001001011000101000: oled_data = 16'b0100100111000111;
				18'b001001011010101000: oled_data = 16'b1011010100110011;
				18'b001001011100101000: oled_data = 16'b1111011101011100;
				18'b001001011110101000: oled_data = 16'b1110111100011011;
				18'b001001100000101000: oled_data = 16'b1110111100011010;
				18'b001001100010101000: oled_data = 16'b1110111100011010;
				18'b001001100100101000: oled_data = 16'b1110111100011010;
				18'b001001100110101000: oled_data = 16'b1110111100011010;
				18'b001001101000101000: oled_data = 16'b1110111100011010;
				18'b001001101010101000: oled_data = 16'b1110111100011010;
				18'b001001101100101000: oled_data = 16'b1110111100011010;
				18'b001001101110101000: oled_data = 16'b1110111100011010;
				18'b001001110000101000: oled_data = 16'b1101111010011000;
				18'b001001110010101000: oled_data = 16'b1110011011111010;
				18'b001001110100101000: oled_data = 16'b1110111100111011;
				18'b001001110110101000: oled_data = 16'b1101111001111000;
				18'b001001111000101000: oled_data = 16'b1101010101110101;
				18'b001001111010101000: oled_data = 16'b1101010101010101;
				18'b001001111100101000: oled_data = 16'b1101110100010100;
				18'b001001111110101000: oled_data = 16'b1100101111001111;
				18'b001010000000101000: oled_data = 16'b1010101000001000;
				18'b001010000010101000: oled_data = 16'b1011101011101011;
				18'b001010000100101000: oled_data = 16'b1110110011110011;
				18'b001010000110101000: oled_data = 16'b1100101101101110;
				18'b001010001000101000: oled_data = 16'b1011001000101001;
				18'b001010001010101000: oled_data = 16'b1011001001001001;
				18'b001010001100101000: oled_data = 16'b1011001001001001;
				18'b001010001110101000: oled_data = 16'b1011001000101001;
				18'b001010010000101000: oled_data = 16'b1011001101101110;
				18'b001010010010101000: oled_data = 16'b1100011011111011;
				18'b001010010100101000: oled_data = 16'b1011111011111011;
				18'b001010010110101000: oled_data = 16'b1011111011111011;
				18'b001010011000101000: oled_data = 16'b1011111011111100;
				18'b001010011010101000: oled_data = 16'b1100011100111100;
				18'b001010011100101000: oled_data = 16'b1011110101010101;
				18'b001010011110101000: oled_data = 16'b1010101000001000;
				18'b001010100000101000: oled_data = 16'b1010101000001000;
				18'b001010100010101000: oled_data = 16'b1010001000001000;
				18'b001010100100101000: oled_data = 16'b1010101000001000;
				18'b001010100110101000: oled_data = 16'b1010101000001000;
				18'b001000011000101001: oled_data = 16'b1101110011010101;
				18'b001000011010101001: oled_data = 16'b1101110011010101;
				18'b001000011100101001: oled_data = 16'b1101110011010101;
				18'b001000011110101001: oled_data = 16'b1101110011010101;
				18'b001000100000101001: oled_data = 16'b1101010001110100;
				18'b001000100010101001: oled_data = 16'b1100110001010011;
				18'b001000100100101001: oled_data = 16'b1011001101110000;
				18'b001000100110101001: oled_data = 16'b1100010001010011;
				18'b001000101000101001: oled_data = 16'b1101010010010101;
				18'b001000101010101001: oled_data = 16'b1100010000110010;
				18'b001000101100101001: oled_data = 16'b1101110011110110;
				18'b001000101110101001: oled_data = 16'b1101110011010101;
				18'b001000110000101001: oled_data = 16'b1101110011010101;
				18'b001000110010101001: oled_data = 16'b1101110011010101;
				18'b001000110100101001: oled_data = 16'b1101110011010101;
				18'b001000110110101001: oled_data = 16'b1101110011010110;
				18'b001000111000101001: oled_data = 16'b1101110010010101;
				18'b001000111010101001: oled_data = 16'b1101010011110101;
				18'b001000111100101001: oled_data = 16'b1110111011111010;
				18'b001000111110101001: oled_data = 16'b1110011100011010;
				18'b001001000000101001: oled_data = 16'b1110111100011010;
				18'b001001000010101001: oled_data = 16'b1110111100011010;
				18'b001001000100101001: oled_data = 16'b1110111100011010;
				18'b001001000110101001: oled_data = 16'b1110111100011010;
				18'b001001001000101001: oled_data = 16'b1110111100011010;
				18'b001001001010101001: oled_data = 16'b1110111100011010;
				18'b001001001100101001: oled_data = 16'b1110111100011010;
				18'b001001001110101001: oled_data = 16'b1110111100011010;
				18'b001001010000101001: oled_data = 16'b1110111100111010;
				18'b001001010010101001: oled_data = 16'b1110011100011010;
				18'b001001010100101001: oled_data = 16'b0111001100101100;
				18'b001001010110101001: oled_data = 16'b0011000100100100;
				18'b001001011000101001: oled_data = 16'b1001010001010000;
				18'b001001011010101001: oled_data = 16'b1110111100111011;
				18'b001001011100101001: oled_data = 16'b1110111100011010;
				18'b001001011110101001: oled_data = 16'b1110111100011010;
				18'b001001100000101001: oled_data = 16'b1110111100011010;
				18'b001001100010101001: oled_data = 16'b1110111100011010;
				18'b001001100100101001: oled_data = 16'b1110111100011010;
				18'b001001100110101001: oled_data = 16'b1110111100011010;
				18'b001001101000101001: oled_data = 16'b1110111100011010;
				18'b001001101010101001: oled_data = 16'b1110111100011010;
				18'b001001101100101001: oled_data = 16'b1110111100011010;
				18'b001001101110101001: oled_data = 16'b1101111010111001;
				18'b001001110000101001: oled_data = 16'b1110011011011001;
				18'b001001110010101001: oled_data = 16'b1110111100111011;
				18'b001001110100101001: oled_data = 16'b1101111010011000;
				18'b001001110110101001: oled_data = 16'b1101010111010110;
				18'b001001111000101001: oled_data = 16'b1110111010111001;
				18'b001001111010101001: oled_data = 16'b1110111011011001;
				18'b001001111100101001: oled_data = 16'b1101110101010100;
				18'b001001111110101001: oled_data = 16'b1100101110001110;
				18'b001010000000101001: oled_data = 16'b1011001000001000;
				18'b001010000010101001: oled_data = 16'b1100101110101110;
				18'b001010000100101001: oled_data = 16'b1110010011010010;
				18'b001010000110101001: oled_data = 16'b1011101010001010;
				18'b001010001000101001: oled_data = 16'b1011001001001001;
				18'b001010001010101001: oled_data = 16'b1011001001001001;
				18'b001010001100101001: oled_data = 16'b1011001001001001;
				18'b001010001110101001: oled_data = 16'b1011001000101001;
				18'b001010010000101001: oled_data = 16'b1011110011010011;
				18'b001010010010101001: oled_data = 16'b1011111100011100;
				18'b001010010100101001: oled_data = 16'b1011111011111011;
				18'b001010010110101001: oled_data = 16'b1011111011111011;
				18'b001010011000101001: oled_data = 16'b1011111011111100;
				18'b001010011010101001: oled_data = 16'b1100111100111101;
				18'b001010011100101001: oled_data = 16'b1100011010011001;
				18'b001010011110101001: oled_data = 16'b1011001011001011;
				18'b001010100000101001: oled_data = 16'b1010101000101000;
				18'b001010100010101001: oled_data = 16'b1010101000101000;
				18'b001010100100101001: oled_data = 16'b1010101000001000;
				18'b001010100110101001: oled_data = 16'b1010101000001000;
				18'b001000011000101010: oled_data = 16'b1101110011010101;
				18'b001000011010101010: oled_data = 16'b1101110011010101;
				18'b001000011100101010: oled_data = 16'b1101110011010101;
				18'b001000011110101010: oled_data = 16'b1101110010110101;
				18'b001000100000101010: oled_data = 16'b1101010001110100;
				18'b001000100010101010: oled_data = 16'b1100001111010010;
				18'b001000100100101010: oled_data = 16'b1011001101110001;
				18'b001000100110101010: oled_data = 16'b1101010001110100;
				18'b001000101000101010: oled_data = 16'b1101010010010100;
				18'b001000101010101010: oled_data = 16'b1011110001010010;
				18'b001000101100101010: oled_data = 16'b1101110011010110;
				18'b001000101110101010: oled_data = 16'b1101110011010110;
				18'b001000110000101010: oled_data = 16'b1101110011010101;
				18'b001000110010101010: oled_data = 16'b1101110011010101;
				18'b001000110100101010: oled_data = 16'b1101110011010101;
				18'b001000110110101010: oled_data = 16'b1101110011010110;
				18'b001000111000101010: oled_data = 16'b1101010010010100;
				18'b001000111010101010: oled_data = 16'b1101010101010110;
				18'b001000111100101010: oled_data = 16'b1110011100011010;
				18'b001000111110101010: oled_data = 16'b1110111100011010;
				18'b001001000000101010: oled_data = 16'b1110111100011010;
				18'b001001000010101010: oled_data = 16'b1110111100011010;
				18'b001001000100101010: oled_data = 16'b1110111100011010;
				18'b001001000110101010: oled_data = 16'b1110111100011010;
				18'b001001001000101010: oled_data = 16'b1110111100011010;
				18'b001001001010101010: oled_data = 16'b1110111100011010;
				18'b001001001100101010: oled_data = 16'b1110111100011010;
				18'b001001001110101010: oled_data = 16'b1110111100011010;
				18'b001001010000101010: oled_data = 16'b1110111100111011;
				18'b001001010010101010: oled_data = 16'b1000001111101111;
				18'b001001010100101010: oled_data = 16'b0011000100100100;
				18'b001001010110101010: oled_data = 16'b0111001100101100;
				18'b001001011000101010: oled_data = 16'b1110011100011011;
				18'b001001011010101010: oled_data = 16'b1110111100011011;
				18'b001001011100101010: oled_data = 16'b1110111100011010;
				18'b001001011110101010: oled_data = 16'b1110111100011010;
				18'b001001100000101010: oled_data = 16'b1110111100011010;
				18'b001001100010101010: oled_data = 16'b1110111100011010;
				18'b001001100100101010: oled_data = 16'b1110111100011010;
				18'b001001100110101010: oled_data = 16'b1110111100011010;
				18'b001001101000101010: oled_data = 16'b1110111100011010;
				18'b001001101010101010: oled_data = 16'b1110111100011010;
				18'b001001101100101010: oled_data = 16'b1110111100011010;
				18'b001001101110101010: oled_data = 16'b1110011011111010;
				18'b001001110000101010: oled_data = 16'b1110111100111010;
				18'b001001110010101010: oled_data = 16'b1101111010011000;
				18'b001001110100101010: oled_data = 16'b1101011000110111;
				18'b001001110110101010: oled_data = 16'b1110111011011010;
				18'b001001111000101010: oled_data = 16'b1110111100011011;
				18'b001001111010101010: oled_data = 16'b1110011011011010;
				18'b001001111100101010: oled_data = 16'b1101010100110100;
				18'b001001111110101010: oled_data = 16'b1100001101001101;
				18'b001010000000101010: oled_data = 16'b1010101000101000;
				18'b001010000010101010: oled_data = 16'b1101010000110000;
				18'b001010000100101010: oled_data = 16'b1101010000010000;
				18'b001010000110101010: oled_data = 16'b1011001001001001;
				18'b001010001000101010: oled_data = 16'b1011101001001001;
				18'b001010001010101010: oled_data = 16'b1011001001001001;
				18'b001010001100101010: oled_data = 16'b1011001001001001;
				18'b001010001110101010: oled_data = 16'b1011001001001001;
				18'b001010010000101010: oled_data = 16'b1100010111010111;
				18'b001010010010101010: oled_data = 16'b1011111100011100;
				18'b001010010100101010: oled_data = 16'b1011111011111011;
				18'b001010010110101010: oled_data = 16'b1011111011111011;
				18'b001010011000101010: oled_data = 16'b1011111011111011;
				18'b001010011010101010: oled_data = 16'b1100111100011100;
				18'b001010011100101010: oled_data = 16'b1011111100011011;
				18'b001010011110101010: oled_data = 16'b1011001111001111;
				18'b001010100000101010: oled_data = 16'b1010101000001000;
				18'b001010100010101010: oled_data = 16'b1010101000101000;
				18'b001010100100101010: oled_data = 16'b1010101000001000;
				18'b001010100110101010: oled_data = 16'b1010101000001000;
				18'b001000011000101011: oled_data = 16'b1101110011010101;
				18'b001000011010101011: oled_data = 16'b1101110011010101;
				18'b001000011100101011: oled_data = 16'b1101110011010101;
				18'b001000011110101011: oled_data = 16'b1101110010010101;
				18'b001000100000101011: oled_data = 16'b1100110000110100;
				18'b001000100010101011: oled_data = 16'b1011101110010001;
				18'b001000100100101011: oled_data = 16'b1011001101110001;
				18'b001000100110101011: oled_data = 16'b1101110010010101;
				18'b001000101000101011: oled_data = 16'b1100110001110011;
				18'b001000101010101011: oled_data = 16'b1100010001010011;
				18'b001000101100101011: oled_data = 16'b1101110011010110;
				18'b001000101110101011: oled_data = 16'b1101110011010110;
				18'b001000110000101011: oled_data = 16'b1101110011010101;
				18'b001000110010101011: oled_data = 16'b1101110011010101;
				18'b001000110100101011: oled_data = 16'b1101110011010101;
				18'b001000110110101011: oled_data = 16'b1101110011010110;
				18'b001000111000101011: oled_data = 16'b1101010010010100;
				18'b001000111010101011: oled_data = 16'b1101010110010111;
				18'b001000111100101011: oled_data = 16'b1110111100011010;
				18'b001000111110101011: oled_data = 16'b1110111100011010;
				18'b001001000000101011: oled_data = 16'b1110111100011010;
				18'b001001000010101011: oled_data = 16'b1110111100011010;
				18'b001001000100101011: oled_data = 16'b1110111100011010;
				18'b001001000110101011: oled_data = 16'b1110111100011010;
				18'b001001001000101011: oled_data = 16'b1110111100011010;
				18'b001001001010101011: oled_data = 16'b1110111100011010;
				18'b001001001100101011: oled_data = 16'b1110111100011010;
				18'b001001001110101011: oled_data = 16'b1110111101011011;
				18'b001001010000101011: oled_data = 16'b1001110010110001;
				18'b001001010010101011: oled_data = 16'b0010100100000100;
				18'b001001010100101011: oled_data = 16'b0110001010101011;
				18'b001001010110101011: oled_data = 16'b1101111010111010;
				18'b001001011000101011: oled_data = 16'b1110111100111011;
				18'b001001011010101011: oled_data = 16'b1110011100011011;
				18'b001001011100101011: oled_data = 16'b1110111100011011;
				18'b001001011110101011: oled_data = 16'b1110111100011011;
				18'b001001100000101011: oled_data = 16'b1110111100011011;
				18'b001001100010101011: oled_data = 16'b1110111100011011;
				18'b001001100100101011: oled_data = 16'b1110111100011011;
				18'b001001100110101011: oled_data = 16'b1110111100011011;
				18'b001001101000101011: oled_data = 16'b1110111100011011;
				18'b001001101010101011: oled_data = 16'b1110111100011011;
				18'b001001101100101011: oled_data = 16'b1110111100011011;
				18'b001001101110101011: oled_data = 16'b1110111100111011;
				18'b001001110000101011: oled_data = 16'b1101011000010111;
				18'b001001110010101011: oled_data = 16'b1101111000010111;
				18'b001001110100101011: oled_data = 16'b1110111011111010;
				18'b001001110110101011: oled_data = 16'b1110111100011010;
				18'b001001111000101011: oled_data = 16'b1110111011111010;
				18'b001001111010101011: oled_data = 16'b1110011011011010;
				18'b001001111100101011: oled_data = 16'b1101010101010100;
				18'b001001111110101011: oled_data = 16'b1011101100001101;
				18'b001010000000101011: oled_data = 16'b1011001000101001;
				18'b001010000010101011: oled_data = 16'b1101110001110001;
				18'b001010000100101011: oled_data = 16'b1100101101101110;
				18'b001010000110101011: oled_data = 16'b1011001000101001;
				18'b001010001000101011: oled_data = 16'b1011101001001001;
				18'b001010001010101011: oled_data = 16'b1011001001001001;
				18'b001010001100101011: oled_data = 16'b1011001000101001;
				18'b001010001110101011: oled_data = 16'b1011001010101011;
				18'b001010010000101011: oled_data = 16'b1100011001111010;
				18'b001010010010101011: oled_data = 16'b1011111011111100;
				18'b001010010100101011: oled_data = 16'b1011111011111011;
				18'b001010010110101011: oled_data = 16'b1011111011111011;
				18'b001010011000101011: oled_data = 16'b1011111011111011;
				18'b001010011010101011: oled_data = 16'b1100111100011100;
				18'b001010011100101011: oled_data = 16'b1011111100011100;
				18'b001010011110101011: oled_data = 16'b1011010011010010;
				18'b001010100000101011: oled_data = 16'b1010101000001000;
				18'b001010100010101011: oled_data = 16'b1010101000001000;
				18'b001010100100101011: oled_data = 16'b1010101000001000;
				18'b001010100110101011: oled_data = 16'b1010101000001000;
				18'b001000011000101100: oled_data = 16'b1101110010110101;
				18'b001000011010101100: oled_data = 16'b1101110010110101;
				18'b001000011100101100: oled_data = 16'b1101110011010101;
				18'b001000011110101100: oled_data = 16'b1101010001110100;
				18'b001000100000101100: oled_data = 16'b1100001111110011;
				18'b001000100010101100: oled_data = 16'b1011001101110001;
				18'b001000100100101100: oled_data = 16'b1011001110010001;
				18'b001000100110101100: oled_data = 16'b1101110010110101;
				18'b001000101000101100: oled_data = 16'b1100110000010011;
				18'b001000101010101100: oled_data = 16'b1100010000110011;
				18'b001000101100101100: oled_data = 16'b1101110011010110;
				18'b001000101110101100: oled_data = 16'b1101110011010110;
				18'b001000110000101100: oled_data = 16'b1101110011010101;
				18'b001000110010101100: oled_data = 16'b1101110011010101;
				18'b001000110100101100: oled_data = 16'b1101110011010101;
				18'b001000110110101100: oled_data = 16'b1101110011010101;
				18'b001000111000101100: oled_data = 16'b1100110001110100;
				18'b001000111010101100: oled_data = 16'b1101010111011000;
				18'b001000111100101100: oled_data = 16'b1110111100011010;
				18'b001000111110101100: oled_data = 16'b1110011100011010;
				18'b001001000000101100: oled_data = 16'b1110011100011010;
				18'b001001000010101100: oled_data = 16'b1110011100011010;
				18'b001001000100101100: oled_data = 16'b1110011100011010;
				18'b001001000110101100: oled_data = 16'b1110011100011010;
				18'b001001001000101100: oled_data = 16'b1110011100011010;
				18'b001001001010101100: oled_data = 16'b1110111100011010;
				18'b001001001100101100: oled_data = 16'b1110111101011011;
				18'b001001001110101100: oled_data = 16'b1010110100010011;
				18'b001001010000101100: oled_data = 16'b0011000101000100;
				18'b001001010010101100: oled_data = 16'b0101001001001001;
				18'b001001010100101100: oled_data = 16'b1101111001111001;
				18'b001001010110101100: oled_data = 16'b1110111100111011;
				18'b001001011000101100: oled_data = 16'b1110011100011010;
				18'b001001011010101100: oled_data = 16'b1110011100011010;
				18'b001001011100101100: oled_data = 16'b1110011100011010;
				18'b001001011110101100: oled_data = 16'b1110011100011010;
				18'b001001100000101100: oled_data = 16'b1110111100011010;
				18'b001001100010101100: oled_data = 16'b1110111100011010;
				18'b001001100100101100: oled_data = 16'b1110111100011010;
				18'b001001100110101100: oled_data = 16'b1110111100011010;
				18'b001001101000101100: oled_data = 16'b1110111100011010;
				18'b001001101010101100: oled_data = 16'b1110111100111011;
				18'b001001101100101100: oled_data = 16'b1110011011011010;
				18'b001001101110101100: oled_data = 16'b1101010110010110;
				18'b001001110000101100: oled_data = 16'b1101010111110110;
				18'b001001110010101100: oled_data = 16'b1110111011111010;
				18'b001001110100101100: oled_data = 16'b1110111011111010;
				18'b001001110110101100: oled_data = 16'b1110011100011010;
				18'b001001111000101100: oled_data = 16'b1110011011111010;
				18'b001001111010101100: oled_data = 16'b1110111100011010;
				18'b001001111100101100: oled_data = 16'b1101010101110101;
				18'b001001111110101100: oled_data = 16'b1011101011101100;
				18'b001010000000101100: oled_data = 16'b1011001001001010;
				18'b001010000010101100: oled_data = 16'b1101110010010010;
				18'b001010000100101100: oled_data = 16'b1100001011101100;
				18'b001010000110101100: oled_data = 16'b1011001000101001;
				18'b001010001000101100: oled_data = 16'b1011001001001001;
				18'b001010001010101100: oled_data = 16'b1011001001001001;
				18'b001010001100101100: oled_data = 16'b1011001000101001;
				18'b001010001110101100: oled_data = 16'b1011101011101100;
				18'b001010010000101100: oled_data = 16'b1100011010111011;
				18'b001010010010101100: oled_data = 16'b1011111011111100;
				18'b001010010100101100: oled_data = 16'b1011111011111011;
				18'b001010010110101100: oled_data = 16'b1011111011111011;
				18'b001010011000101100: oled_data = 16'b1011111011111011;
				18'b001010011010101100: oled_data = 16'b1011111011111011;
				18'b001010011100101100: oled_data = 16'b1011111100011100;
				18'b001010011110101100: oled_data = 16'b1011110100010100;
				18'b001010100000101100: oled_data = 16'b1010101000001000;
				18'b001010100010101100: oled_data = 16'b1010101000001000;
				18'b001010100100101100: oled_data = 16'b1010101000001000;
				18'b001010100110101100: oled_data = 16'b1010101000001000;
				18'b001000011000101101: oled_data = 16'b1101110010110101;
				18'b001000011010101101: oled_data = 16'b1101110010110101;
				18'b001000011100101101: oled_data = 16'b1101110010110101;
				18'b001000011110101101: oled_data = 16'b1100110001010100;
				18'b001000100000101101: oled_data = 16'b1100001111010010;
				18'b001000100010101101: oled_data = 16'b1011001101110001;
				18'b001000100100101101: oled_data = 16'b1011001110010001;
				18'b001000100110101101: oled_data = 16'b1101110010110101;
				18'b001000101000101101: oled_data = 16'b1100010000010010;
				18'b001000101010101101: oled_data = 16'b1100110000110011;
				18'b001000101100101101: oled_data = 16'b1101110011010110;
				18'b001000101110101101: oled_data = 16'b1101110011010110;
				18'b001000110000101101: oled_data = 16'b1101110011010101;
				18'b001000110010101101: oled_data = 16'b1101110011010101;
				18'b001000110100101101: oled_data = 16'b1101110011010101;
				18'b001000110110101101: oled_data = 16'b1101110011010101;
				18'b001000111000101101: oled_data = 16'b1100110001110100;
				18'b001000111010101101: oled_data = 16'b1101111000011000;
				18'b001000111100101101: oled_data = 16'b1110111100011010;
				18'b001000111110101101: oled_data = 16'b1110011100011010;
				18'b001001000000101101: oled_data = 16'b1110011100011010;
				18'b001001000010101101: oled_data = 16'b1110011100011010;
				18'b001001000100101101: oled_data = 16'b1110011100011010;
				18'b001001000110101101: oled_data = 16'b1110011100011010;
				18'b001001001000101101: oled_data = 16'b1110011100011010;
				18'b001001001010101101: oled_data = 16'b1110111100111010;
				18'b001001001100101101: oled_data = 16'b1100010110010101;
				18'b001001001110101101: oled_data = 16'b0011100101100101;
				18'b001001010000101101: oled_data = 16'b0100101000101000;
				18'b001001010010101101: oled_data = 16'b1101011000111000;
				18'b001001010100101101: oled_data = 16'b1110111100111011;
				18'b001001010110101101: oled_data = 16'b1110011100011010;
				18'b001001011000101101: oled_data = 16'b1110011100011010;
				18'b001001011010101101: oled_data = 16'b1110011100011010;
				18'b001001011100101101: oled_data = 16'b1110011100011010;
				18'b001001011110101101: oled_data = 16'b1110011100011010;
				18'b001001100000101101: oled_data = 16'b1110111100011010;
				18'b001001100010101101: oled_data = 16'b1110111100011010;
				18'b001001100100101101: oled_data = 16'b1110011100011010;
				18'b001001100110101101: oled_data = 16'b1110111100111010;
				18'b001001101000101101: oled_data = 16'b1110111100111011;
				18'b001001101010101101: oled_data = 16'b1101111000110111;
				18'b001001101100101101: oled_data = 16'b1101010100110100;
				18'b001001101110101101: oled_data = 16'b1101110101010101;
				18'b001001110000101101: oled_data = 16'b1110111011011010;
				18'b001001110010101101: oled_data = 16'b1110111100011010;
				18'b001001110100101101: oled_data = 16'b1110111011111010;
				18'b001001110110101101: oled_data = 16'b1110011100011010;
				18'b001001111000101101: oled_data = 16'b1110011100011010;
				18'b001001111010101101: oled_data = 16'b1110111100011010;
				18'b001001111100101101: oled_data = 16'b1101010110110110;
				18'b001001111110101101: oled_data = 16'b1011101011001100;
				18'b001010000000101101: oled_data = 16'b1011001001001010;
				18'b001010000010101101: oled_data = 16'b1101110001110001;
				18'b001010000100101101: oled_data = 16'b1011101010001011;
				18'b001010000110101101: oled_data = 16'b1011001001001001;
				18'b001010001000101101: oled_data = 16'b1011001001001001;
				18'b001010001010101101: oled_data = 16'b1011001001001001;
				18'b001010001100101101: oled_data = 16'b1011001000101001;
				18'b001010001110101101: oled_data = 16'b1011101100001100;
				18'b001010010000101101: oled_data = 16'b1100011010111011;
				18'b001010010010101101: oled_data = 16'b1011111011111100;
				18'b001010010100101101: oled_data = 16'b1011111011111100;
				18'b001010010110101101: oled_data = 16'b1010111010011010;
				18'b001010011000101101: oled_data = 16'b1010011000111001;
				18'b001010011010101101: oled_data = 16'b1011011010011010;
				18'b001010011100101101: oled_data = 16'b1011111100111100;
				18'b001010011110101101: oled_data = 16'b1011110100010100;
				18'b001010100000101101: oled_data = 16'b1010101000001000;
				18'b001010100010101101: oled_data = 16'b1010101000001000;
				18'b001010100100101101: oled_data = 16'b1010101000001000;
				18'b001010100110101101: oled_data = 16'b1010101000001000;
				18'b001000011000101110: oled_data = 16'b1101110010110101;
				18'b001000011010101110: oled_data = 16'b1101110010110101;
				18'b001000011100101110: oled_data = 16'b1101110010110101;
				18'b001000011110101110: oled_data = 16'b1100110000110011;
				18'b001000100000101110: oled_data = 16'b1011101110010001;
				18'b001000100010101110: oled_data = 16'b1011001101110001;
				18'b001000100100101110: oled_data = 16'b1011101110110010;
				18'b001000100110101110: oled_data = 16'b1101110010110101;
				18'b001000101000101110: oled_data = 16'b1100001111110010;
				18'b001000101010101110: oled_data = 16'b1100110000110011;
				18'b001000101100101110: oled_data = 16'b1101110011010110;
				18'b001000101110101110: oled_data = 16'b1101110010110101;
				18'b001000110000101110: oled_data = 16'b1101110010110101;
				18'b001000110010101110: oled_data = 16'b1101110010110101;
				18'b001000110100101110: oled_data = 16'b1101110011010101;
				18'b001000110110101110: oled_data = 16'b1101110011010101;
				18'b001000111000101110: oled_data = 16'b1100110001110011;
				18'b001000111010101110: oled_data = 16'b1101111001011000;
				18'b001000111100101110: oled_data = 16'b1110011100011010;
				18'b001000111110101110: oled_data = 16'b1110011100011010;
				18'b001001000000101110: oled_data = 16'b1110011100011010;
				18'b001001000010101110: oled_data = 16'b1110011100011010;
				18'b001001000100101110: oled_data = 16'b1110011011111010;
				18'b001001000110101110: oled_data = 16'b1110011011111010;
				18'b001001001000101110: oled_data = 16'b1110011100011010;
				18'b001001001010101110: oled_data = 16'b1101111011011001;
				18'b001001001100101110: oled_data = 16'b1100110111010110;
				18'b001001001110101110: oled_data = 16'b1001110010110001;
				18'b001001010000101110: oled_data = 16'b1101011001011000;
				18'b001001010010101110: oled_data = 16'b1110111100111011;
				18'b001001010100101110: oled_data = 16'b1110011100011010;
				18'b001001010110101110: oled_data = 16'b1110011100011010;
				18'b001001011000101110: oled_data = 16'b1110011100011010;
				18'b001001011010101110: oled_data = 16'b1110011100011010;
				18'b001001011100101110: oled_data = 16'b1110011011111010;
				18'b001001011110101110: oled_data = 16'b1110011100011010;
				18'b001001100000101110: oled_data = 16'b1110011100011010;
				18'b001001100010101110: oled_data = 16'b1110111100011010;
				18'b001001100100101110: oled_data = 16'b1110011100011010;
				18'b001001100110101110: oled_data = 16'b1101111001011000;
				18'b001001101000101110: oled_data = 16'b1100010011010011;
				18'b001001101010101110: oled_data = 16'b1100110001110010;
				18'b001001101100101110: oled_data = 16'b1101010011110100;
				18'b001001101110101110: oled_data = 16'b1110010111110111;
				18'b001001110000101110: oled_data = 16'b1110111011111010;
				18'b001001110010101110: oled_data = 16'b1110011011111010;
				18'b001001110100101110: oled_data = 16'b1110111011111010;
				18'b001001110110101110: oled_data = 16'b1110011011111010;
				18'b001001111000101110: oled_data = 16'b1110011011111010;
				18'b001001111010101110: oled_data = 16'b1110111100011010;
				18'b001001111100101110: oled_data = 16'b1101111000110111;
				18'b001001111110101110: oled_data = 16'b1011001011001011;
				18'b001010000000101110: oled_data = 16'b1011001001101010;
				18'b001010000010101110: oled_data = 16'b1101010000110000;
				18'b001010000100101110: oled_data = 16'b1011101001101010;
				18'b001010000110101110: oled_data = 16'b1011001001001001;
				18'b001010001000101110: oled_data = 16'b1011001001001001;
				18'b001010001010101110: oled_data = 16'b1011001001001001;
				18'b001010001100101110: oled_data = 16'b1011001000101001;
				18'b001010001110101110: oled_data = 16'b1011101011001100;
				18'b001010010000101110: oled_data = 16'b1100011010011011;
				18'b001010010010101110: oled_data = 16'b1011111011111100;
				18'b001010010100101110: oled_data = 16'b1011011010011011;
				18'b001010010110101110: oled_data = 16'b1001010111011000;
				18'b001010011000101110: oled_data = 16'b1001010110111000;
				18'b001010011010101110: oled_data = 16'b1010111001011010;
				18'b001010011100101110: oled_data = 16'b1011011011111100;
				18'b001010011110101110: oled_data = 16'b1011010010110010;
				18'b001010100000101110: oled_data = 16'b1010100111101000;
				18'b001010100010101110: oled_data = 16'b1010101000001000;
				18'b001010100100101110: oled_data = 16'b1010101000001000;
				18'b001010100110101110: oled_data = 16'b1010101000001000;
				18'b001000011000101111: oled_data = 16'b1101110010010101;
				18'b001000011010101111: oled_data = 16'b1101110010010101;
				18'b001000011100101111: oled_data = 16'b1101010010010101;
				18'b001000011110101111: oled_data = 16'b1100001111110010;
				18'b001000100000101111: oled_data = 16'b1011001101010000;
				18'b001000100010101111: oled_data = 16'b1011001101010000;
				18'b001000100100101111: oled_data = 16'b1011101110110001;
				18'b001000100110101111: oled_data = 16'b1101110011010101;
				18'b001000101000101111: oled_data = 16'b1100001111010010;
				18'b001000101010101111: oled_data = 16'b1100110000110011;
				18'b001000101100101111: oled_data = 16'b1101110010110110;
				18'b001000101110101111: oled_data = 16'b1101110010110101;
				18'b001000110000101111: oled_data = 16'b1101110010110101;
				18'b001000110010101111: oled_data = 16'b1101110010110101;
				18'b001000110100101111: oled_data = 16'b1101110010110101;
				18'b001000110110101111: oled_data = 16'b1101110010110101;
				18'b001000111000101111: oled_data = 16'b1100110001110011;
				18'b001000111010101111: oled_data = 16'b1101111001111000;
				18'b001000111100101111: oled_data = 16'b1110011100011010;
				18'b001000111110101111: oled_data = 16'b1110011011111010;
				18'b001001000000101111: oled_data = 16'b1110111100111010;
				18'b001001000010101111: oled_data = 16'b1110011100011010;
				18'b001001000100101111: oled_data = 16'b1110011011111010;
				18'b001001000110101111: oled_data = 16'b1110011011111010;
				18'b001001001000101111: oled_data = 16'b1110011011111010;
				18'b001001001010101111: oled_data = 16'b1110011011111010;
				18'b001001001100101111: oled_data = 16'b1110111100011010;
				18'b001001001110101111: oled_data = 16'b1110111100111010;
				18'b001001010000101111: oled_data = 16'b1110011100011010;
				18'b001001010010101111: oled_data = 16'b1110011011111010;
				18'b001001010100101111: oled_data = 16'b1110011011111010;
				18'b001001010110101111: oled_data = 16'b1110011011111010;
				18'b001001011000101111: oled_data = 16'b1110011100011010;
				18'b001001011010101111: oled_data = 16'b1110011100011010;
				18'b001001011100101111: oled_data = 16'b1110111100011010;
				18'b001001011110101111: oled_data = 16'b1110111100011010;
				18'b001001100000101111: oled_data = 16'b1110011011011001;
				18'b001001100010101111: oled_data = 16'b1101010111110110;
				18'b001001100100101111: oled_data = 16'b1011110010010010;
				18'b001001100110101111: oled_data = 16'b1011001111001111;
				18'b001001101000101111: oled_data = 16'b1100110001010010;
				18'b001001101010101111: oled_data = 16'b1101110011110100;
				18'b001001101100101111: oled_data = 16'b1101010011110100;
				18'b001001101110101111: oled_data = 16'b1110111001011000;
				18'b001001110000101111: oled_data = 16'b1110011010111001;
				18'b001001110010101111: oled_data = 16'b1110011011111010;
				18'b001001110100101111: oled_data = 16'b1110011011111010;
				18'b001001110110101111: oled_data = 16'b1110011011111010;
				18'b001001111000101111: oled_data = 16'b1110011011111010;
				18'b001001111010101111: oled_data = 16'b1110011100011010;
				18'b001001111100101111: oled_data = 16'b1110011011111001;
				18'b001001111110101111: oled_data = 16'b1010101100101100;
				18'b001010000000101111: oled_data = 16'b1011001001101010;
				18'b001010000010101111: oled_data = 16'b1100101111101111;
				18'b001010000100101111: oled_data = 16'b1011001001001001;
				18'b001010000110101111: oled_data = 16'b1011001001001001;
				18'b001010001000101111: oled_data = 16'b1011001001101001;
				18'b001010001010101111: oled_data = 16'b1011001001001001;
				18'b001010001100101111: oled_data = 16'b1011001000101001;
				18'b001010001110101111: oled_data = 16'b1011001001001010;
				18'b001010010000101111: oled_data = 16'b1100011000011000;
				18'b001010010010101111: oled_data = 16'b1011111100011100;
				18'b001010010100101111: oled_data = 16'b1010011000111001;
				18'b001010010110101111: oled_data = 16'b1001010111011000;
				18'b001010011000101111: oled_data = 16'b1001010111011000;
				18'b001010011010101111: oled_data = 16'b1001110111011000;
				18'b001010011100101111: oled_data = 16'b1010111001111010;
				18'b001010011110101111: oled_data = 16'b1011001110101111;
				18'b001010100000101111: oled_data = 16'b1010100111101000;
				18'b001010100010101111: oled_data = 16'b1010100111101000;
				18'b001010100100101111: oled_data = 16'b1010101000001000;
				18'b001010100110101111: oled_data = 16'b1010100111101000;
				18'b001000011000110000: oled_data = 16'b1101010010010100;
				18'b001000011010110000: oled_data = 16'b1101010010010100;
				18'b001000011100110000: oled_data = 16'b1101010001010100;
				18'b001000011110110000: oled_data = 16'b1011101110010001;
				18'b001000100000110000: oled_data = 16'b1010101100110000;
				18'b001000100010110000: oled_data = 16'b1010101100110000;
				18'b001000100100110000: oled_data = 16'b1011101110110010;
				18'b001000100110110000: oled_data = 16'b1101110011010101;
				18'b001000101000110000: oled_data = 16'b1011101110110001;
				18'b001000101010110000: oled_data = 16'b1100110000010011;
				18'b001000101100110000: oled_data = 16'b1101110010110110;
				18'b001000101110110000: oled_data = 16'b1101110010010101;
				18'b001000110000110000: oled_data = 16'b1101010001110100;
				18'b001000110010110000: oled_data = 16'b1101010001110100;
				18'b001000110100110000: oled_data = 16'b1101110010110101;
				18'b001000110110110000: oled_data = 16'b1101110010110101;
				18'b001000111000110000: oled_data = 16'b1100110001110011;
				18'b001000111010110000: oled_data = 16'b1110011010011001;
				18'b001000111100110000: oled_data = 16'b1100010101110101;
				18'b001000111110110000: oled_data = 16'b1010110001010001;
				18'b001001000000110000: oled_data = 16'b1100110101110101;
				18'b001001000010110000: oled_data = 16'b1101111001111000;
				18'b001001000100110000: oled_data = 16'b1110011011011010;
				18'b001001000110110000: oled_data = 16'b1110011011111010;
				18'b001001001000110000: oled_data = 16'b1110011100011010;
				18'b001001001010110000: oled_data = 16'b1110011100011010;
				18'b001001001100110000: oled_data = 16'b1110011100011010;
				18'b001001001110110000: oled_data = 16'b1110011100011010;
				18'b001001010000110000: oled_data = 16'b1110111100011010;
				18'b001001010010110000: oled_data = 16'b1110011100011010;
				18'b001001010100110000: oled_data = 16'b1110011100011010;
				18'b001001010110110000: oled_data = 16'b1110011100011010;
				18'b001001011000110000: oled_data = 16'b1110011011111010;
				18'b001001011010110000: oled_data = 16'b1101111010011000;
				18'b001001011100110000: oled_data = 16'b1101010111010110;
				18'b001001011110110000: oled_data = 16'b1100010011110011;
				18'b001001100000110000: oled_data = 16'b1011110000010000;
				18'b001001100010110000: oled_data = 16'b1011001110001111;
				18'b001001100100110000: oled_data = 16'b1011001110001111;
				18'b001001100110110000: oled_data = 16'b1100110001010010;
				18'b001001101000110000: oled_data = 16'b1101110100010101;
				18'b001001101010110000: oled_data = 16'b1100110010110011;
				18'b001001101100110000: oled_data = 16'b1101010011110100;
				18'b001001101110110000: oled_data = 16'b1101010101110101;
				18'b001001110000110000: oled_data = 16'b1101111001111000;
				18'b001001110010110000: oled_data = 16'b1110011011111010;
				18'b001001110100110000: oled_data = 16'b1110011011111010;
				18'b001001110110110000: oled_data = 16'b1110011011111010;
				18'b001001111000110000: oled_data = 16'b1110011011111010;
				18'b001001111010110000: oled_data = 16'b1110011011111010;
				18'b001001111100110000: oled_data = 16'b1110011011111001;
				18'b001001111110110000: oled_data = 16'b1011001110101110;
				18'b001010000000110000: oled_data = 16'b1011001001101010;
				18'b001010000010110000: oled_data = 16'b1100101110001110;
				18'b001010000100110000: oled_data = 16'b1011001000101001;
				18'b001010000110110000: oled_data = 16'b1011001000101001;
				18'b001010001000110000: oled_data = 16'b1100101101101101;
				18'b001010001010110000: oled_data = 16'b1011101001101010;
				18'b001010001100110000: oled_data = 16'b1011001000101001;
				18'b001010001110110000: oled_data = 16'b1011001000001000;
				18'b001010010000110000: oled_data = 16'b1011110001010001;
				18'b001010010010110000: oled_data = 16'b1011111100111100;
				18'b001010010100110000: oled_data = 16'b1001111000111001;
				18'b001010010110110000: oled_data = 16'b1001010110110111;
				18'b001010011000110000: oled_data = 16'b1001010111010111;
				18'b001010011010110000: oled_data = 16'b1001010111111000;
				18'b001010011100110000: oled_data = 16'b1011010101110110;
				18'b001010011110110000: oled_data = 16'b1010101001001001;
				18'b001010100000110000: oled_data = 16'b1010000111101000;
				18'b001010100010110000: oled_data = 16'b1010000111000111;
				18'b001010100100110000: oled_data = 16'b1001100111000111;
				18'b001010100110110000: oled_data = 16'b1001100111000111;
				18'b001000011000110001: oled_data = 16'b1101010001110100;
				18'b001000011010110001: oled_data = 16'b1101010001110100;
				18'b001000011100110001: oled_data = 16'b1100010000010011;
				18'b001000011110110001: oled_data = 16'b1011001101010000;
				18'b001000100000110001: oled_data = 16'b1010101100001111;
				18'b001000100010110001: oled_data = 16'b1010101100001111;
				18'b001000100100110001: oled_data = 16'b1011101110110010;
				18'b001000100110110001: oled_data = 16'b1101110010110101;
				18'b001000101000110001: oled_data = 16'b1011101110110001;
				18'b001000101010110001: oled_data = 16'b1100001111110010;
				18'b001000101100110001: oled_data = 16'b1101110010110110;
				18'b001000101110110001: oled_data = 16'b1101110010010101;
				18'b001000110000110001: oled_data = 16'b1101010001010100;
				18'b001000110010110001: oled_data = 16'b1100110000110011;
				18'b001000110100110001: oled_data = 16'b1101010010010101;
				18'b001000110110110001: oled_data = 16'b1101010010010100;
				18'b001000111000110001: oled_data = 16'b1100010000010010;
				18'b001000111010110001: oled_data = 16'b1011010000010001;
				18'b001000111100110001: oled_data = 16'b1011001110001111;
				18'b001000111110110001: oled_data = 16'b1011101110010000;
				18'b001001000000110001: oled_data = 16'b1011001101101111;
				18'b001001000010110001: oled_data = 16'b1011001110001111;
				18'b001001000100110001: oled_data = 16'b1011010000010000;
				18'b001001000110110001: oled_data = 16'b1011010010110010;
				18'b001001001000110001: oled_data = 16'b1011110101110100;
				18'b001001001010110001: oled_data = 16'b1100111000110111;
				18'b001001001100110001: oled_data = 16'b1101011001010111;
				18'b001001001110110001: oled_data = 16'b1101011000010111;
				18'b001001010000110001: oled_data = 16'b1100010110110101;
				18'b001001010010110001: oled_data = 16'b1100010101010101;
				18'b001001010100110001: oled_data = 16'b1100010100110100;
				18'b001001010110110001: oled_data = 16'b1011110011010010;
				18'b001001011000110001: oled_data = 16'b1011010001110001;
				18'b001001011010110001: oled_data = 16'b1010101111001111;
				18'b001001011100110001: oled_data = 16'b1011001110001111;
				18'b001001011110110001: oled_data = 16'b1011101110001111;
				18'b001001100000110001: oled_data = 16'b1011101110110000;
				18'b001001100010110001: oled_data = 16'b1011101110110000;
				18'b001001100100110001: oled_data = 16'b1100110001110010;
				18'b001001100110110001: oled_data = 16'b1110010100010101;
				18'b001001101000110001: oled_data = 16'b1101010010110011;
				18'b001001101010110001: oled_data = 16'b1101010011010011;
				18'b001001101100110001: oled_data = 16'b1100110010110011;
				18'b001001101110110001: oled_data = 16'b1100110100010100;
				18'b001001110000110001: oled_data = 16'b1101111001111000;
				18'b001001110010110001: oled_data = 16'b1110011011011001;
				18'b001001110100110001: oled_data = 16'b1110011011111010;
				18'b001001110110110001: oled_data = 16'b1110011011111010;
				18'b001001111000110001: oled_data = 16'b1110011011111010;
				18'b001001111010110001: oled_data = 16'b1110011011011001;
				18'b001001111100110001: oled_data = 16'b1110011011111010;
				18'b001001111110110001: oled_data = 16'b1011101111001111;
				18'b001010000000110001: oled_data = 16'b1011001001001001;
				18'b001010000010110001: oled_data = 16'b1100001101001101;
				18'b001010000100110001: oled_data = 16'b1011001000101001;
				18'b001010000110110001: oled_data = 16'b1011001001001001;
				18'b001010001000110001: oled_data = 16'b1100101101101101;
				18'b001010001010110001: oled_data = 16'b1011001001001001;
				18'b001010001100110001: oled_data = 16'b1011001000101000;
				18'b001010001110110001: oled_data = 16'b1011001000101001;
				18'b001010010000110001: oled_data = 16'b1001100111101000;
				18'b001010010010110001: oled_data = 16'b1010110011110011;
				18'b001010010100110001: oled_data = 16'b1011011001111010;
				18'b001010010110110001: oled_data = 16'b1001010111111000;
				18'b001010011000110001: oled_data = 16'b1001010111011000;
				18'b001010011010110001: oled_data = 16'b1010010101110110;
				18'b001010011100110001: oled_data = 16'b1001001001101001;
				18'b001010011110110001: oled_data = 16'b1000100101100101;
				18'b001010100000110001: oled_data = 16'b1010000111000111;
				18'b001010100010110001: oled_data = 16'b1010100111101000;
				18'b001010100100110001: oled_data = 16'b1010000111100111;
				18'b001010100110110001: oled_data = 16'b1010000111000111;
				18'b001000011000110010: oled_data = 16'b1101010000110011;
				18'b001000011010110010: oled_data = 16'b1101010001010100;
				18'b001000011100110010: oled_data = 16'b1011101111010010;
				18'b001000011110110010: oled_data = 16'b1010101100001111;
				18'b001000100000110010: oled_data = 16'b1010101011101111;
				18'b001000100010110010: oled_data = 16'b1010001011101111;
				18'b001000100100110010: oled_data = 16'b1011101110110010;
				18'b001000100110110010: oled_data = 16'b1101010010010101;
				18'b001000101000110010: oled_data = 16'b1011101110110001;
				18'b001000101010110010: oled_data = 16'b1011101110110001;
				18'b001000101100110010: oled_data = 16'b1101110010010101;
				18'b001000101110110010: oled_data = 16'b1101010001110100;
				18'b001000110000110010: oled_data = 16'b1101010001010100;
				18'b001000110010110010: oled_data = 16'b1100110000010011;
				18'b001000110100110010: oled_data = 16'b1101010001110100;
				18'b001000110110110010: oled_data = 16'b1101010001110100;
				18'b001000111000110010: oled_data = 16'b1011101110110001;
				18'b001000111010110010: oled_data = 16'b1010101101001111;
				18'b001000111100110010: oled_data = 16'b1011101110110000;
				18'b001000111110110010: oled_data = 16'b1011101110110000;
				18'b001001000000110010: oled_data = 16'b1011101110010000;
				18'b001001000010110010: oled_data = 16'b1011001110001111;
				18'b001001000100110010: oled_data = 16'b1010101101001110;
				18'b001001000110110010: oled_data = 16'b1011110001010001;
				18'b001001001000110010: oled_data = 16'b1101010111110110;
				18'b001001001010110010: oled_data = 16'b1101111010011000;
				18'b001001001100110010: oled_data = 16'b1101111010111001;
				18'b001001001110110010: oled_data = 16'b1110011010011001;
				18'b001001010000110010: oled_data = 16'b1101010111010110;
				18'b001001010010110010: oled_data = 16'b1100010001110010;
				18'b001001010100110010: oled_data = 16'b1011101110101111;
				18'b001001010110110010: oled_data = 16'b1011001110001111;
				18'b001001011000110010: oled_data = 16'b1011101110001111;
				18'b001001011010110010: oled_data = 16'b1011101111010000;
				18'b001001011100110010: oled_data = 16'b1011101110110000;
				18'b001001011110110010: oled_data = 16'b1011101111010000;
				18'b001001100000110010: oled_data = 16'b1100010000010001;
				18'b001001100010110010: oled_data = 16'b1100110001110010;
				18'b001001100100110010: oled_data = 16'b1101110011110100;
				18'b001001100110110010: oled_data = 16'b1101010011010100;
				18'b001001101000110010: oled_data = 16'b1100110010010011;
				18'b001001101010110010: oled_data = 16'b1101110100010101;
				18'b001001101100110010: oled_data = 16'b1100110010110011;
				18'b001001101110110010: oled_data = 16'b1100010011010011;
				18'b001001110000110010: oled_data = 16'b1101010111010110;
				18'b001001110010110010: oled_data = 16'b1110011010111001;
				18'b001001110100110010: oled_data = 16'b1110011011011001;
				18'b001001110110110010: oled_data = 16'b1110011011011001;
				18'b001001111000110010: oled_data = 16'b1101111010011000;
				18'b001001111010110010: oled_data = 16'b1101011001111000;
				18'b001001111100110010: oled_data = 16'b1110011010011001;
				18'b001001111110110010: oled_data = 16'b1011001101101101;
				18'b001010000000110010: oled_data = 16'b1011001001001001;
				18'b001010000010110010: oled_data = 16'b1100001100101100;
				18'b001010000100110010: oled_data = 16'b1011001000101001;
				18'b001010000110110010: oled_data = 16'b1011001001001001;
				18'b001010001000110010: oled_data = 16'b1011101010101010;
				18'b001010001010110010: oled_data = 16'b1011001000101000;
				18'b001010001100110010: oled_data = 16'b1011001000001000;
				18'b001010001110110010: oled_data = 16'b1011001000101000;
				18'b001010010000110010: oled_data = 16'b1001000110100111;
				18'b001010010010110010: oled_data = 16'b1001000111000111;
				18'b001010010100110010: oled_data = 16'b1011001100101101;
				18'b001010010110110010: oled_data = 16'b1010101110101111;
				18'b001010011000110010: oled_data = 16'b1010101100101101;
				18'b001010011010110010: oled_data = 16'b1010001001001001;
				18'b001010011100110010: oled_data = 16'b1010000111000111;
				18'b001010011110110010: oled_data = 16'b1010000111000111;
				18'b001010100000110010: oled_data = 16'b1010000111000111;
				18'b001010100010110010: oled_data = 16'b1010000111000111;
				18'b001010100100110010: oled_data = 16'b1010000111000111;
				18'b001010100110110010: oled_data = 16'b1010000111000111;
				18'b001000011000110011: oled_data = 16'b1100110000010011;
				18'b001000011010110011: oled_data = 16'b1101010000110011;
				18'b001000011100110011: oled_data = 16'b1011001101010000;
				18'b001000011110110011: oled_data = 16'b1010001011001110;
				18'b001000100000110011: oled_data = 16'b1010001011101111;
				18'b001000100010110011: oled_data = 16'b1010001011101111;
				18'b001000100100110011: oled_data = 16'b1011101110110010;
				18'b001000100110110011: oled_data = 16'b1101010001110100;
				18'b001000101000110011: oled_data = 16'b1011001110010001;
				18'b001000101010110011: oled_data = 16'b1011001101010000;
				18'b001000101100110011: oled_data = 16'b1101010001010100;
				18'b001000101110110011: oled_data = 16'b1101010000110100;
				18'b001000110000110011: oled_data = 16'b1100110000110011;
				18'b001000110010110011: oled_data = 16'b1100001111110010;
				18'b001000110100110011: oled_data = 16'b1101010000110011;
				18'b001000110110110011: oled_data = 16'b1101010001010100;
				18'b001000111000110011: oled_data = 16'b1011101110010000;
				18'b001000111010110011: oled_data = 16'b1010001011101101;
				18'b001000111100110011: oled_data = 16'b1010101100001110;
				18'b001000111110110011: oled_data = 16'b1011001101001110;
				18'b001001000000110011: oled_data = 16'b1011001110001111;
				18'b001001000010110011: oled_data = 16'b1011001101101111;
				18'b001001000100110011: oled_data = 16'b1011110010010010;
				18'b001001000110110011: oled_data = 16'b1101111010011001;
				18'b001001001000110011: oled_data = 16'b1110011011011001;
				18'b001001001010110011: oled_data = 16'b1110011010111001;
				18'b001001001100110011: oled_data = 16'b1110011011011001;
				18'b001001001110110011: oled_data = 16'b1110011011011001;
				18'b001001010000110011: oled_data = 16'b1110011011011010;
				18'b001001010010110011: oled_data = 16'b1101111010011001;
				18'b001001010100110011: oled_data = 16'b1011110011110011;
				18'b001001010110110011: oled_data = 16'b1011001111110000;
				18'b001001011000110011: oled_data = 16'b1011001110001111;
				18'b001001011010110011: oled_data = 16'b1011001110001111;
				18'b001001011100110011: oled_data = 16'b1011101111010000;
				18'b001001011110110011: oled_data = 16'b1100110001110010;
				18'b001001100000110011: oled_data = 16'b1101110011010100;
				18'b001001100010110011: oled_data = 16'b1100110010110011;
				18'b001001100100110011: oled_data = 16'b1101010010010011;
				18'b001001100110110011: oled_data = 16'b1100110010010010;
				18'b001001101000110011: oled_data = 16'b1101010011010100;
				18'b001001101010110011: oled_data = 16'b1101010011110100;
				18'b001001101100110011: oled_data = 16'b1100110010110011;
				18'b001001101110110011: oled_data = 16'b1100110010110011;
				18'b001001110000110011: oled_data = 16'b1100110011110100;
				18'b001001110010110011: oled_data = 16'b1100010101010100;
				18'b001001110100110011: oled_data = 16'b1101010111010110;
				18'b001001110110110011: oled_data = 16'b1100110111110110;
				18'b001001111000110011: oled_data = 16'b1101011000110111;
				18'b001001111010110011: oled_data = 16'b1101110111110111;
				18'b001001111100110011: oled_data = 16'b1101010100110101;
				18'b001001111110110011: oled_data = 16'b1011001011101100;
				18'b001010000000110011: oled_data = 16'b1011001001001001;
				18'b001010000010110011: oled_data = 16'b1011101100001100;
				18'b001010000100110011: oled_data = 16'b1010101000001000;
				18'b001010000110110011: oled_data = 16'b1011001000001000;
				18'b001010001000110011: oled_data = 16'b1011001000001000;
				18'b001010001010110011: oled_data = 16'b1011001000001000;
				18'b001010001100110011: oled_data = 16'b1010101000001000;
				18'b001010001110110011: oled_data = 16'b1010101000001000;
				18'b001010010000110011: oled_data = 16'b1001000110000110;
				18'b001010010010110011: oled_data = 16'b1010000111001000;
				18'b001010010100110011: oled_data = 16'b1010100111100111;
				18'b001010010110110011: oled_data = 16'b1010100111000111;
				18'b001010011000110011: oled_data = 16'b1010000111000111;
				18'b001010011010110011: oled_data = 16'b1010000111100111;
				18'b001010011100110011: oled_data = 16'b1010000111100111;
				18'b001010011110110011: oled_data = 16'b1010000111000111;
				18'b001010100000110011: oled_data = 16'b1010000111000111;
				18'b001010100010110011: oled_data = 16'b1001100111000111;
				18'b001010100100110011: oled_data = 16'b1001100111000111;
				18'b001010100110110011: oled_data = 16'b1001100111000111;
				18'b001000011000110100: oled_data = 16'b1100101111110011;
				18'b001000011010110100: oled_data = 16'b1100101111110011;
				18'b001000011100110100: oled_data = 16'b1011001100001111;
				18'b001000011110110100: oled_data = 16'b1010001010101110;
				18'b001000100000110100: oled_data = 16'b1001101010101110;
				18'b001000100010110100: oled_data = 16'b1001101010101110;
				18'b001000100100110100: oled_data = 16'b1011101110010001;
				18'b001000100110110100: oled_data = 16'b1101010001010100;
				18'b001000101000110100: oled_data = 16'b1011001101110000;
				18'b001000101010110100: oled_data = 16'b1010001100001111;
				18'b001000101100110100: oled_data = 16'b1100110000110100;
				18'b001000101110110100: oled_data = 16'b1100110000010011;
				18'b001000110000110100: oled_data = 16'b1100110000010011;
				18'b001000110010110100: oled_data = 16'b1100001111010010;
				18'b001000110100110100: oled_data = 16'b1100110000010011;
				18'b001000110110110100: oled_data = 16'b1101010000110011;
				18'b001000111000110100: oled_data = 16'b1011001110010000;
				18'b001000111010110100: oled_data = 16'b1010101100101110;
				18'b001000111100110100: oled_data = 16'b1010101100101110;
				18'b001000111110110100: oled_data = 16'b1010101100101110;
				18'b001001000000110100: oled_data = 16'b1010101011101101;
				18'b001001000010110100: oled_data = 16'b1010101111001111;
				18'b001001000100110100: oled_data = 16'b1101011001011000;
				18'b001001000110110100: oled_data = 16'b1101111010111001;
				18'b001001001000110100: oled_data = 16'b1101111010111001;
				18'b001001001010110100: oled_data = 16'b1101111010111001;
				18'b001001001100110100: oled_data = 16'b1101111010111001;
				18'b001001001110110100: oled_data = 16'b1101111010111001;
				18'b001001010000110100: oled_data = 16'b1101111010111001;
				18'b001001010010110100: oled_data = 16'b1101011010011000;
				18'b001001010100110100: oled_data = 16'b1101011000010111;
				18'b001001010110110100: oled_data = 16'b1011110001110001;
				18'b001001011000110100: oled_data = 16'b1011001110001111;
				18'b001001011010110100: oled_data = 16'b1011101111010000;
				18'b001001011100110100: oled_data = 16'b1100010000110001;
				18'b001001011110110100: oled_data = 16'b1100110001110010;
				18'b001001100000110100: oled_data = 16'b1100110010010011;
				18'b001001100010110100: oled_data = 16'b1011110000010001;
				18'b001001100100110100: oled_data = 16'b1100110001010010;
				18'b001001100110110100: oled_data = 16'b1101010011010100;
				18'b001001101000110100: oled_data = 16'b1101010011010100;
				18'b001001101010110100: oled_data = 16'b1101010011010100;
				18'b001001101100110100: oled_data = 16'b1101010010110100;
				18'b001001101110110100: oled_data = 16'b1100110010010011;
				18'b001001110000110100: oled_data = 16'b1100110010010011;
				18'b001001110010110100: oled_data = 16'b1011110001110010;
				18'b001001110100110100: oled_data = 16'b1100010010110011;
				18'b001001110110110100: oled_data = 16'b1101010101010101;
				18'b001001111000110100: oled_data = 16'b1100110100110100;
				18'b001001111010110100: oled_data = 16'b1100110010110011;
				18'b001001111100110100: oled_data = 16'b1101010010110100;
				18'b001001111110110100: oled_data = 16'b1010101011101100;
				18'b001010000000110100: oled_data = 16'b1011001000101000;
				18'b001010000010110100: oled_data = 16'b1011001011001011;
				18'b001010000100110100: oled_data = 16'b1010101000001000;
				18'b001010000110110100: oled_data = 16'b1010101000001000;
				18'b001010001000110100: oled_data = 16'b1010101000001000;
				18'b001010001010110100: oled_data = 16'b1010101000001000;
				18'b001010001100110100: oled_data = 16'b1010101000001000;
				18'b001010001110110100: oled_data = 16'b1010101000001000;
				18'b001010010000110100: oled_data = 16'b1000100110000110;
				18'b001010010010110100: oled_data = 16'b1010000111101000;
				18'b001010010100110100: oled_data = 16'b1010100111101000;
				18'b001010010110110100: oled_data = 16'b1010000111101000;
				18'b001010011000110100: oled_data = 16'b1010000111001000;
				18'b001010011010110100: oled_data = 16'b1010000111000111;
				18'b001010011100110100: oled_data = 16'b1010000111000111;
				18'b001010011110110100: oled_data = 16'b1010000111000111;
				18'b001010100000110100: oled_data = 16'b1010000111000111;
				18'b001010100010110100: oled_data = 16'b1001100111000111;
				18'b001010100100110100: oled_data = 16'b1001100110100111;
				18'b001010100110110100: oled_data = 16'b1001100110100111;
				18'b001000011000110101: oled_data = 16'b1100001111010010;
				18'b001000011010110101: oled_data = 16'b1100001111010010;
				18'b001000011100110101: oled_data = 16'b1010101011001110;
				18'b001000011110110101: oled_data = 16'b1001101010101101;
				18'b001000100000110101: oled_data = 16'b1001101010001101;
				18'b001000100010110101: oled_data = 16'b1001101010001101;
				18'b001000100100110101: oled_data = 16'b1011001101110001;
				18'b001000100110110101: oled_data = 16'b1100110000110011;
				18'b001000101000110101: oled_data = 16'b1011001101010000;
				18'b001000101010110101: oled_data = 16'b1001101010101110;
				18'b001000101100110101: oled_data = 16'b1100001111110010;
				18'b001000101110110101: oled_data = 16'b1100010000010011;
				18'b001000110000110101: oled_data = 16'b1100110000010011;
				18'b001000110010110101: oled_data = 16'b1100001111010010;
				18'b001000110100110101: oled_data = 16'b1100001111010010;
				18'b001000110110110101: oled_data = 16'b1101010000010011;
				18'b001000111000110101: oled_data = 16'b1011001110010000;
				18'b001000111010110101: oled_data = 16'b1011101111110001;
				18'b001000111100110101: oled_data = 16'b1011101111110001;
				18'b001000111110110101: oled_data = 16'b1011101110010000;
				18'b001001000000110101: oled_data = 16'b1010101101101111;
				18'b001001000010110101: oled_data = 16'b1100110110010101;
				18'b001001000100110101: oled_data = 16'b1101111010011001;
				18'b001001000110110101: oled_data = 16'b1101111010011000;
				18'b001001001000110101: oled_data = 16'b1101111010011000;
				18'b001001001010110101: oled_data = 16'b1101111010011000;
				18'b001001001100110101: oled_data = 16'b1101111010011000;
				18'b001001001110110101: oled_data = 16'b1101111010011000;
				18'b001001010000110101: oled_data = 16'b1101111010011000;
				18'b001001010010110101: oled_data = 16'b1101111010011000;
				18'b001001010100110101: oled_data = 16'b1101011000110111;
				18'b001001010110110101: oled_data = 16'b1100110100010100;
				18'b001001011000110101: oled_data = 16'b1101010010110011;
				18'b001001011010110101: oled_data = 16'b1101010010110011;
				18'b001001011100110101: oled_data = 16'b1101010010110011;
				18'b001001011110110101: oled_data = 16'b1100110010010010;
				18'b001001100000110101: oled_data = 16'b1100010001110010;
				18'b001001100010110101: oled_data = 16'b1011110000010001;
				18'b001001100100110101: oled_data = 16'b1101010010110011;
				18'b001001100110110101: oled_data = 16'b1101010010110011;
				18'b001001101000110101: oled_data = 16'b1101010010110011;
				18'b001001101010110101: oled_data = 16'b1101010010110011;
				18'b001001101100110101: oled_data = 16'b1101010010110011;
				18'b001001101110110101: oled_data = 16'b1100010001010010;
				18'b001001110000110101: oled_data = 16'b1100110001110010;
				18'b001001110010110101: oled_data = 16'b1100110010010011;
				18'b001001110100110101: oled_data = 16'b1100110010010011;
				18'b001001110110110101: oled_data = 16'b1101010010110011;
				18'b001001111000110101: oled_data = 16'b1101010010110011;
				18'b001001111010110101: oled_data = 16'b1100110010010011;
				18'b001001111100110101: oled_data = 16'b1100010000110010;
				18'b001001111110110101: oled_data = 16'b1010101010101011;
				18'b001010000000110101: oled_data = 16'b1011001000001000;
				18'b001010000010110101: oled_data = 16'b1011001010101010;
				18'b001010000100110101: oled_data = 16'b1010101000001000;
				18'b001010000110110101: oled_data = 16'b1010101000001000;
				18'b001010001000110101: oled_data = 16'b1010101000001000;
				18'b001010001010110101: oled_data = 16'b1010101000001000;
				18'b001010001100110101: oled_data = 16'b1010100111101000;
				18'b001010001110110101: oled_data = 16'b1010000111101000;
				18'b001010010000110101: oled_data = 16'b1000100110000110;
				18'b001010010010110101: oled_data = 16'b1010000111101000;
				18'b001010010100110101: oled_data = 16'b1010000111101000;
				18'b001010010110110101: oled_data = 16'b1010000111000111;
				18'b001010011000110101: oled_data = 16'b1001100111000111;
				18'b001010011010110101: oled_data = 16'b1001100111000111;
				18'b001010011100110101: oled_data = 16'b1001100111000111;
				18'b001010011110110101: oled_data = 16'b1001100110100111;
				18'b001010100000110101: oled_data = 16'b1001100110100111;
				18'b001010100010110101: oled_data = 16'b1001100110100111;
				18'b001010100100110101: oled_data = 16'b1001100110100111;
				18'b001010100110110101: oled_data = 16'b1001100110100111;
				18'b001000011000110110: oled_data = 16'b1100001110110010;
				18'b001000011010110110: oled_data = 16'b1100001111010010;
				18'b001000011100110110: oled_data = 16'b1010001010101110;
				18'b001000011110110110: oled_data = 16'b1001101010001101;
				18'b001000100000110110: oled_data = 16'b1001001010001101;
				18'b001000100010110110: oled_data = 16'b1001001010001101;
				18'b001000100100110110: oled_data = 16'b1011001101010000;
				18'b001000100110110110: oled_data = 16'b1100001111110011;
				18'b001000101000110110: oled_data = 16'b1011001101110000;
				18'b001000101010110110: oled_data = 16'b1001001010001101;
				18'b001000101100110110: oled_data = 16'b1011101110110001;
				18'b001000101110110110: oled_data = 16'b1100001111110010;
				18'b001000110000110110: oled_data = 16'b1100001111110010;
				18'b001000110010110110: oled_data = 16'b1100001111010010;
				18'b001000110100110110: oled_data = 16'b1011101101110001;
				18'b001000110110110110: oled_data = 16'b1100101111110010;
				18'b001000111000110110: oled_data = 16'b1011101110010000;
				18'b001000111010110110: oled_data = 16'b1100010000010010;
				18'b001000111100110110: oled_data = 16'b1100110001110011;
				18'b001000111110110110: oled_data = 16'b1100010000110010;
				18'b001001000000110110: oled_data = 16'b1011010001110010;
				18'b001001000010110110: oled_data = 16'b1101011001011000;
				18'b001001000100110110: oled_data = 16'b1101011001111000;
				18'b001001000110110110: oled_data = 16'b1101011001111000;
				18'b001001001000110110: oled_data = 16'b1101011001111000;
				18'b001001001010110110: oled_data = 16'b1101011001111000;
				18'b001001001100110110: oled_data = 16'b1101011001111000;
				18'b001001001110110110: oled_data = 16'b1101011001111000;
				18'b001001010000110110: oled_data = 16'b1101011001111000;
				18'b001001010010110110: oled_data = 16'b1101011001111000;
				18'b001001010100110110: oled_data = 16'b1101111001111000;
				18'b001001010110110110: oled_data = 16'b1100110101010101;
				18'b001001011000110110: oled_data = 16'b1100110010010011;
				18'b001001011010110110: oled_data = 16'b1101010010010011;
				18'b001001011100110110: oled_data = 16'b1100110010010011;
				18'b001001011110110110: oled_data = 16'b1100110010010010;
				18'b001001100000110110: oled_data = 16'b1100110010010010;
				18'b001001100010110110: oled_data = 16'b1100010000110001;
				18'b001001100100110110: oled_data = 16'b1100110010010011;
				18'b001001100110110110: oled_data = 16'b1100110010010011;
				18'b001001101000110110: oled_data = 16'b1100110010010011;
				18'b001001101010110110: oled_data = 16'b1100110010010011;
				18'b001001101100110110: oled_data = 16'b1100110010010011;
				18'b001001101110110110: oled_data = 16'b1100110010010011;
				18'b001001110000110110: oled_data = 16'b1100010000110001;
				18'b001001110010110110: oled_data = 16'b1011001111110000;
				18'b001001110100110110: oled_data = 16'b1011110000110001;
				18'b001001110110110110: oled_data = 16'b1100010001010010;
				18'b001001111000110110: oled_data = 16'b1100010000110001;
				18'b001001111010110110: oled_data = 16'b1100010000010001;
				18'b001001111100110110: oled_data = 16'b1100010001010011;
				18'b001001111110110110: oled_data = 16'b1010101011001100;
				18'b001010000000110110: oled_data = 16'b1010101000001000;
				18'b001010000010110110: oled_data = 16'b1010101001101001;
				18'b001010000100110110: oled_data = 16'b1010100111101000;
				18'b001010000110110110: oled_data = 16'b1010100111101000;
				18'b001010001000110110: oled_data = 16'b1010100111101000;
				18'b001010001010110110: oled_data = 16'b1010000111101000;
				18'b001010001100110110: oled_data = 16'b1010100111100111;
				18'b001010001110110110: oled_data = 16'b1001100111000111;
				18'b001010010000110110: oled_data = 16'b1000100110000110;
				18'b001010010010110110: oled_data = 16'b1010000111000111;
				18'b001010010100110110: oled_data = 16'b1010000111000111;
				18'b001010010110110110: oled_data = 16'b1001100111000111;
				18'b001010011000110110: oled_data = 16'b1001000110100110;
				18'b001010011010110110: oled_data = 16'b1001100110100111;
				18'b001010011100110110: oled_data = 16'b1001100110100111;
				18'b001010011110110110: oled_data = 16'b1001100110100111;
				18'b001010100000110110: oled_data = 16'b1001100110100110;
				18'b001010100010110110: oled_data = 16'b1001100110100110;
				18'b001010100100110110: oled_data = 16'b1001000110100110;
				18'b001010100110110110: oled_data = 16'b1001000110000110;
				18'b001000011000110111: oled_data = 16'b1100001110110001;
				18'b001000011010110111: oled_data = 16'b1100001110110001;
				18'b001000011100110111: oled_data = 16'b1001101010101101;
				18'b001000011110110111: oled_data = 16'b1001001010001100;
				18'b001000100000110111: oled_data = 16'b1001001010001101;
				18'b001000100010110111: oled_data = 16'b1001001010001101;
				18'b001000100100110111: oled_data = 16'b1010101100110000;
				18'b001000100110110111: oled_data = 16'b1100001111010010;
				18'b001000101000110111: oled_data = 16'b1011001101110000;
				18'b001000101010110111: oled_data = 16'b1001001010001101;
				18'b001000101100110111: oled_data = 16'b1010101101110000;
				18'b001000101110110111: oled_data = 16'b1100001111110010;
				18'b001000110000110111: oled_data = 16'b1100001111010010;
				18'b001000110010110111: oled_data = 16'b1011101110110001;
				18'b001000110100110111: oled_data = 16'b1011001101010000;
				18'b001000110110110111: oled_data = 16'b1100001111010010;
				18'b001000111000110111: oled_data = 16'b1011101110110001;
				18'b001000111010110111: oled_data = 16'b1100010000010010;
				18'b001000111100110111: oled_data = 16'b1100110001010011;
				18'b001000111110110111: oled_data = 16'b1100010000010001;
				18'b001001000000110111: oled_data = 16'b1100010011010011;
				18'b001001000010110111: oled_data = 16'b1101011000110111;
				18'b001001000100110111: oled_data = 16'b1101011001011000;
				18'b001001000110110111: oled_data = 16'b1101011001011000;
				18'b001001001000110111: oled_data = 16'b1101011001011000;
				18'b001001001010110111: oled_data = 16'b1101011001010111;
				18'b001001001100110111: oled_data = 16'b1101011001010111;
				18'b001001001110110111: oled_data = 16'b1101011001010111;
				18'b001001010000110111: oled_data = 16'b1101011001010111;
				18'b001001010010110111: oled_data = 16'b1101011001010111;
				18'b001001010100110111: oled_data = 16'b1101011000110111;
				18'b001001010110110111: oled_data = 16'b1100110011110011;
				18'b001001011000110111: oled_data = 16'b1100110010010010;
				18'b001001011010110111: oled_data = 16'b1100110001110010;
				18'b001001011100110111: oled_data = 16'b1100110001110010;
				18'b001001011110110111: oled_data = 16'b1100110001110010;
				18'b001001100000110111: oled_data = 16'b1100110001110010;
				18'b001001100010110111: oled_data = 16'b1100010000010001;
				18'b001001100100110111: oled_data = 16'b1100110001110010;
				18'b001001100110110111: oled_data = 16'b1100110001110010;
				18'b001001101000110111: oled_data = 16'b1100110001110011;
				18'b001001101010110111: oled_data = 16'b1100110001010011;
				18'b001001101100110111: oled_data = 16'b1100110001110011;
				18'b001001101110110111: oled_data = 16'b1100110001110011;
				18'b001001110000110111: oled_data = 16'b1011001111110001;
				18'b001001110010110111: oled_data = 16'b0110000111001000;
				18'b001001110100110111: oled_data = 16'b1010101111010000;
				18'b001001110110110111: oled_data = 16'b1011110000010001;
				18'b001001111000110111: oled_data = 16'b1011110000010001;
				18'b001001111010110111: oled_data = 16'b1100110001110010;
				18'b001001111100110111: oled_data = 16'b1100110001110011;
				18'b001001111110110111: oled_data = 16'b1010101011001011;
				18'b001010000000110111: oled_data = 16'b1010101000001000;
				18'b001010000010110111: oled_data = 16'b1010001000101000;
				18'b001010000100110111: oled_data = 16'b1010100111101000;
				18'b001010000110110111: oled_data = 16'b1010100111100111;
				18'b001010001000110111: oled_data = 16'b1010000111100111;
				18'b001010001010110111: oled_data = 16'b1010000111100111;
				18'b001010001100110111: oled_data = 16'b1010000111000111;
				18'b001010001110110111: oled_data = 16'b1001100110100111;
				18'b001010010000110111: oled_data = 16'b1000100110000111;
				18'b001010010010110111: oled_data = 16'b1010000111001000;
				18'b001010010100110111: oled_data = 16'b1010000111000111;
				18'b001010010110110111: oled_data = 16'b1001100111000111;
				18'b001010011000110111: oled_data = 16'b1001000110100110;
				18'b001010011010110111: oled_data = 16'b1001100110100111;
				18'b001010011100110111: oled_data = 16'b1001100110100111;
				18'b001010011110110111: oled_data = 16'b1001100110100110;
				18'b001010100000110111: oled_data = 16'b1001100110000110;
				18'b001010100010110111: oled_data = 16'b1001000110000110;
				18'b001010100100110111: oled_data = 16'b1001000110000110;
				18'b001010100110110111: oled_data = 16'b1001000110000110;
				18'b001100011000001000: oled_data = 16'b1001101111101011;
				18'b001100011010001000: oled_data = 16'b1010010000001011;
				18'b001100011100001000: oled_data = 16'b1010010000101011;
				18'b001100011110001000: oled_data = 16'b1010110000101011;
				18'b001100100000001000: oled_data = 16'b1010110001001101;
				18'b001100100010001000: oled_data = 16'b1110011000111001;
				18'b001100100100001000: oled_data = 16'b1110010101010111;
				18'b001100100110001000: oled_data = 16'b1101110011010101;
				18'b001100101000001000: oled_data = 16'b1101110011010101;
				18'b001100101010001000: oled_data = 16'b1101110011010101;
				18'b001100101100001000: oled_data = 16'b1101110011010101;
				18'b001100101110001000: oled_data = 16'b1101110011010101;
				18'b001100110000001000: oled_data = 16'b1101110011010101;
				18'b001100110010001000: oled_data = 16'b1101110011010101;
				18'b001100110100001000: oled_data = 16'b1101110011010101;
				18'b001100110110001000: oled_data = 16'b1101110011010101;
				18'b001100111000001000: oled_data = 16'b1101110011010101;
				18'b001100111010001000: oled_data = 16'b1101110011010101;
				18'b001100111100001000: oled_data = 16'b1101110011010101;
				18'b001100111110001000: oled_data = 16'b1101110011010101;
				18'b001101000000001000: oled_data = 16'b1101110011010101;
				18'b001101000010001000: oled_data = 16'b1101110011010101;
				18'b001101000100001000: oled_data = 16'b1101110011010101;
				18'b001101000110001000: oled_data = 16'b1101110011010101;
				18'b001101001000001000: oled_data = 16'b1101110011010101;
				18'b001101001010001000: oled_data = 16'b1101110011010101;
				18'b001101001100001000: oled_data = 16'b1101110011010101;
				18'b001101001110001000: oled_data = 16'b1101110011010101;
				18'b001101010000001000: oled_data = 16'b1101110011010101;
				18'b001101010010001000: oled_data = 16'b1101110011010101;
				18'b001101010100001000: oled_data = 16'b1101110011010101;
				18'b001101010110001000: oled_data = 16'b1101110011010101;
				18'b001101011000001000: oled_data = 16'b1101110011010101;
				18'b001101011010001000: oled_data = 16'b1101110011010101;
				18'b001101011100001000: oled_data = 16'b1101110011010101;
				18'b001101011110001000: oled_data = 16'b1101110011010101;
				18'b001101100000001000: oled_data = 16'b1101110011010101;
				18'b001101100010001000: oled_data = 16'b1101110011010101;
				18'b001101100100001000: oled_data = 16'b1101110011010101;
				18'b001101100110001000: oled_data = 16'b1101110011010101;
				18'b001101101000001000: oled_data = 16'b1101110011010101;
				18'b001101101010001000: oled_data = 16'b1101110011010101;
				18'b001101101100001000: oled_data = 16'b1101110011010101;
				18'b001101101110001000: oled_data = 16'b1101110011010101;
				18'b001101110000001000: oled_data = 16'b1101110010110101;
				18'b001101110010001000: oled_data = 16'b1101110011010110;
				18'b001101110100001000: oled_data = 16'b1111011000111010;
				18'b001101110110001000: oled_data = 16'b1100010111010111;
				18'b001101111000001000: oled_data = 16'b1010010100110100;
				18'b001101111010001000: oled_data = 16'b1010010100110100;
				18'b001101111100001000: oled_data = 16'b0101101011101011;
				18'b001101111110001000: oled_data = 16'b0100001000000111;
				18'b001110000000001000: oled_data = 16'b0100001000001000;
				18'b001110000010001000: oled_data = 16'b0100001000001000;
				18'b001110000100001000: oled_data = 16'b0100001000000111;
				18'b001110000110001000: oled_data = 16'b0011100110100110;
				18'b001110001000001000: oled_data = 16'b0101000111100101;
				18'b001110001010001000: oled_data = 16'b0110001001100110;
				18'b001110001100001000: oled_data = 16'b0111001011000110;
				18'b001110001110001000: oled_data = 16'b0111101100000111;
				18'b001110010000001000: oled_data = 16'b0111101100000111;
				18'b001110010010001000: oled_data = 16'b0111101100000111;
				18'b001110010100001000: oled_data = 16'b0111001100001000;
				18'b001110010110001000: oled_data = 16'b0111001011101000;
				18'b001110011000001000: oled_data = 16'b0110101011101000;
				18'b001110011010001000: oled_data = 16'b0110001011001000;
				18'b001110011100001000: oled_data = 16'b0110001010101000;
				18'b001110011110001000: oled_data = 16'b0101101010001000;
				18'b001110100000001000: oled_data = 16'b0101101010001000;
				18'b001110100010001000: oled_data = 16'b0101001001101000;
				18'b001110100100001000: oled_data = 16'b0101001001001000;
				18'b001110100110001000: oled_data = 16'b0101001001101000;
				18'b001100011000001001: oled_data = 16'b1011010001101011;
				18'b001100011010001001: oled_data = 16'b1011010001101011;
				18'b001100011100001001: oled_data = 16'b1011010001001011;
				18'b001100011110001001: oled_data = 16'b1010110000101011;
				18'b001100100000001001: oled_data = 16'b1101010101110100;
				18'b001100100010001001: oled_data = 16'b1110010110011000;
				18'b001100100100001001: oled_data = 16'b1101110011010101;
				18'b001100100110001001: oled_data = 16'b1101110011010101;
				18'b001100101000001001: oled_data = 16'b1101110011010101;
				18'b001100101010001001: oled_data = 16'b1101110011010101;
				18'b001100101100001001: oled_data = 16'b1101110011010101;
				18'b001100101110001001: oled_data = 16'b1101110011010101;
				18'b001100110000001001: oled_data = 16'b1101110011010101;
				18'b001100110010001001: oled_data = 16'b1101110011010101;
				18'b001100110100001001: oled_data = 16'b1101110011010101;
				18'b001100110110001001: oled_data = 16'b1101110011010101;
				18'b001100111000001001: oled_data = 16'b1101110011010101;
				18'b001100111010001001: oled_data = 16'b1101110011010101;
				18'b001100111100001001: oled_data = 16'b1101110011010101;
				18'b001100111110001001: oled_data = 16'b1101110011010101;
				18'b001101000000001001: oled_data = 16'b1101110011010101;
				18'b001101000010001001: oled_data = 16'b1101110011010101;
				18'b001101000100001001: oled_data = 16'b1101110011010101;
				18'b001101000110001001: oled_data = 16'b1101110011010101;
				18'b001101001000001001: oled_data = 16'b1101110011010101;
				18'b001101001010001001: oled_data = 16'b1101110011010101;
				18'b001101001100001001: oled_data = 16'b1101110011010101;
				18'b001101001110001001: oled_data = 16'b1101110011010101;
				18'b001101010000001001: oled_data = 16'b1101110011010101;
				18'b001101010010001001: oled_data = 16'b1101110011010101;
				18'b001101010100001001: oled_data = 16'b1101110011010101;
				18'b001101010110001001: oled_data = 16'b1101110011010101;
				18'b001101011000001001: oled_data = 16'b1101110011010101;
				18'b001101011010001001: oled_data = 16'b1101110011010101;
				18'b001101011100001001: oled_data = 16'b1101110011010101;
				18'b001101011110001001: oled_data = 16'b1101110011010101;
				18'b001101100000001001: oled_data = 16'b1101110011010101;
				18'b001101100010001001: oled_data = 16'b1101110011010101;
				18'b001101100100001001: oled_data = 16'b1101110011010101;
				18'b001101100110001001: oled_data = 16'b1101110011010101;
				18'b001101101000001001: oled_data = 16'b1101110011010101;
				18'b001101101010001001: oled_data = 16'b1101110011010101;
				18'b001101101100001001: oled_data = 16'b1101110011010101;
				18'b001101101110001001: oled_data = 16'b1101110011010101;
				18'b001101110000001001: oled_data = 16'b1101110011010101;
				18'b001101110010001001: oled_data = 16'b1101110010110101;
				18'b001101110100001001: oled_data = 16'b1110010100110111;
				18'b001101110110001001: oled_data = 16'b1110111010011010;
				18'b001101111000001001: oled_data = 16'b1010010011110011;
				18'b001101111010001001: oled_data = 16'b0110101110001101;
				18'b001101111100001001: oled_data = 16'b0100101001101001;
				18'b001101111110001001: oled_data = 16'b0100001000000111;
				18'b001110000000001001: oled_data = 16'b0100001000001000;
				18'b001110000010001001: oled_data = 16'b0100001000001000;
				18'b001110000100001001: oled_data = 16'b0100001000000111;
				18'b001110000110001001: oled_data = 16'b0011100110100101;
				18'b001110001000001001: oled_data = 16'b0100100111000100;
				18'b001110001010001001: oled_data = 16'b0101101001000101;
				18'b001110001100001001: oled_data = 16'b0111001011000111;
				18'b001110001110001001: oled_data = 16'b0111101100000111;
				18'b001110010000001001: oled_data = 16'b1000001100000111;
				18'b001110010010001001: oled_data = 16'b1000001100101000;
				18'b001110010100001001: oled_data = 16'b1000001100101000;
				18'b001110010110001001: oled_data = 16'b1000101101001000;
				18'b001110011000001001: oled_data = 16'b1000101101101000;
				18'b001110011010001001: oled_data = 16'b1000101101101000;
				18'b001110011100001001: oled_data = 16'b1000101101101000;
				18'b001110011110001001: oled_data = 16'b1000101110001001;
				18'b001110100000001001: oled_data = 16'b1000101110001010;
				18'b001110100010001001: oled_data = 16'b0101101010101000;
				18'b001110100100001001: oled_data = 16'b0011101000000111;
				18'b001110100110001001: oled_data = 16'b0100001000101000;
				18'b001100011000001010: oled_data = 16'b1011010001101011;
				18'b001100011010001010: oled_data = 16'b1011010001101011;
				18'b001100011100001010: oled_data = 16'b1010110000101011;
				18'b001100011110001010: oled_data = 16'b1100010011010001;
				18'b001100100000001010: oled_data = 16'b1101110101010111;
				18'b001100100010001010: oled_data = 16'b1101010010110101;
				18'b001100100100001010: oled_data = 16'b1101110011010101;
				18'b001100100110001010: oled_data = 16'b1101110011010101;
				18'b001100101000001010: oled_data = 16'b1101110011010101;
				18'b001100101010001010: oled_data = 16'b1101110011010101;
				18'b001100101100001010: oled_data = 16'b1101110011010101;
				18'b001100101110001010: oled_data = 16'b1101110011010101;
				18'b001100110000001010: oled_data = 16'b1101110011010101;
				18'b001100110010001010: oled_data = 16'b1101110011010101;
				18'b001100110100001010: oled_data = 16'b1101110011010101;
				18'b001100110110001010: oled_data = 16'b1101110011010101;
				18'b001100111000001010: oled_data = 16'b1101110011010101;
				18'b001100111010001010: oled_data = 16'b1101110011010101;
				18'b001100111100001010: oled_data = 16'b1101110011010101;
				18'b001100111110001010: oled_data = 16'b1101110011010101;
				18'b001101000000001010: oled_data = 16'b1101110011010101;
				18'b001101000010001010: oled_data = 16'b1101110011010101;
				18'b001101000100001010: oled_data = 16'b1101110011010101;
				18'b001101000110001010: oled_data = 16'b1101110011010101;
				18'b001101001000001010: oled_data = 16'b1101110011010101;
				18'b001101001010001010: oled_data = 16'b1101110011010101;
				18'b001101001100001010: oled_data = 16'b1101110011010101;
				18'b001101001110001010: oled_data = 16'b1101110011010101;
				18'b001101010000001010: oled_data = 16'b1101110011010101;
				18'b001101010010001010: oled_data = 16'b1101110011010101;
				18'b001101010100001010: oled_data = 16'b1101110011010101;
				18'b001101010110001010: oled_data = 16'b1101110011010101;
				18'b001101011000001010: oled_data = 16'b1101110011010101;
				18'b001101011010001010: oled_data = 16'b1101110011010101;
				18'b001101011100001010: oled_data = 16'b1101110011010101;
				18'b001101011110001010: oled_data = 16'b1101110011010101;
				18'b001101100000001010: oled_data = 16'b1101110011010101;
				18'b001101100010001010: oled_data = 16'b1101110011010101;
				18'b001101100100001010: oled_data = 16'b1101110011010101;
				18'b001101100110001010: oled_data = 16'b1101110011010101;
				18'b001101101000001010: oled_data = 16'b1101110011010110;
				18'b001101101010001010: oled_data = 16'b1101110011010110;
				18'b001101101100001010: oled_data = 16'b1110010011010110;
				18'b001101101110001010: oled_data = 16'b1101110011010101;
				18'b001101110000001010: oled_data = 16'b1101110011010101;
				18'b001101110010001010: oled_data = 16'b1101110011010101;
				18'b001101110100001010: oled_data = 16'b1101110011010101;
				18'b001101110110001010: oled_data = 16'b1110110110111000;
				18'b001101111000001010: oled_data = 16'b1100110111010111;
				18'b001101111010001010: oled_data = 16'b0100101001001001;
				18'b001101111100001010: oled_data = 16'b0100001000000111;
				18'b001101111110001010: oled_data = 16'b0100001000000111;
				18'b001110000000001010: oled_data = 16'b0100001000000111;
				18'b001110000010001010: oled_data = 16'b0100001000000111;
				18'b001110000100001010: oled_data = 16'b0100001000100111;
				18'b001110000110001010: oled_data = 16'b0011000110000101;
				18'b001110001000001010: oled_data = 16'b0010100100100100;
				18'b001110001010001010: oled_data = 16'b0011000101100101;
				18'b001110001100001010: oled_data = 16'b0100000111000110;
				18'b001110001110001010: oled_data = 16'b0101001000000110;
				18'b001110010000001010: oled_data = 16'b0101101001100111;
				18'b001110010010001010: oled_data = 16'b0110101010101000;
				18'b001110010100001010: oled_data = 16'b0111101011101000;
				18'b001110010110001010: oled_data = 16'b1000001100100111;
				18'b001110011000001010: oled_data = 16'b1000101101001000;
				18'b001110011010001010: oled_data = 16'b1000101101101000;
				18'b001110011100001010: oled_data = 16'b1000101110001000;
				18'b001110011110001010: oled_data = 16'b1000101110001000;
				18'b001110100000001010: oled_data = 16'b1000101110001001;
				18'b001110100010001010: oled_data = 16'b0111001011101001;
				18'b001110100100001010: oled_data = 16'b1001001101001101;
				18'b001110100110001010: oled_data = 16'b1011110000010001;
				18'b001100011000001011: oled_data = 16'b1001001111001010;
				18'b001100011010001011: oled_data = 16'b1000101101101001;
				18'b001100011100001011: oled_data = 16'b1001001111001011;
				18'b001100011110001011: oled_data = 16'b1101010100110110;
				18'b001100100000001011: oled_data = 16'b1100110010010100;
				18'b001100100010001011: oled_data = 16'b1101110011010101;
				18'b001100100100001011: oled_data = 16'b1101110011010110;
				18'b001100100110001011: oled_data = 16'b1101110010110101;
				18'b001100101000001011: oled_data = 16'b1101010010010100;
				18'b001100101010001011: oled_data = 16'b1101110011010110;
				18'b001100101100001011: oled_data = 16'b1101110011010101;
				18'b001100101110001011: oled_data = 16'b1101110011010101;
				18'b001100110000001011: oled_data = 16'b1101110011010101;
				18'b001100110010001011: oled_data = 16'b1101110011010101;
				18'b001100110100001011: oled_data = 16'b1101110011010101;
				18'b001100110110001011: oled_data = 16'b1101110011010101;
				18'b001100111000001011: oled_data = 16'b1101110011010101;
				18'b001100111010001011: oled_data = 16'b1101110011010101;
				18'b001100111100001011: oled_data = 16'b1101110011010101;
				18'b001100111110001011: oled_data = 16'b1101110011010101;
				18'b001101000000001011: oled_data = 16'b1101110011010101;
				18'b001101000010001011: oled_data = 16'b1101110011010101;
				18'b001101000100001011: oled_data = 16'b1101110011010101;
				18'b001101000110001011: oled_data = 16'b1101110011010101;
				18'b001101001000001011: oled_data = 16'b1101110011010101;
				18'b001101001010001011: oled_data = 16'b1101110011010101;
				18'b001101001100001011: oled_data = 16'b1101110011010101;
				18'b001101001110001011: oled_data = 16'b1101110011010101;
				18'b001101010000001011: oled_data = 16'b1101110011010101;
				18'b001101010010001011: oled_data = 16'b1101110011010101;
				18'b001101010100001011: oled_data = 16'b1101110011010101;
				18'b001101010110001011: oled_data = 16'b1101110011010101;
				18'b001101011000001011: oled_data = 16'b1101110011010101;
				18'b001101011010001011: oled_data = 16'b1101110011010101;
				18'b001101011100001011: oled_data = 16'b1101110011010101;
				18'b001101011110001011: oled_data = 16'b1101110011010101;
				18'b001101100000001011: oled_data = 16'b1101110011010101;
				18'b001101100010001011: oled_data = 16'b1101110011010101;
				18'b001101100100001011: oled_data = 16'b1101110011010101;
				18'b001101100110001011: oled_data = 16'b1110010011010110;
				18'b001101101000001011: oled_data = 16'b1110010011110110;
				18'b001101101010001011: oled_data = 16'b1110010011110110;
				18'b001101101100001011: oled_data = 16'b1110010011010110;
				18'b001101101110001011: oled_data = 16'b1101110011010101;
				18'b001101110000001011: oled_data = 16'b1101110011010101;
				18'b001101110010001011: oled_data = 16'b1101110011010101;
				18'b001101110100001011: oled_data = 16'b1101110011010101;
				18'b001101110110001011: oled_data = 16'b1101110011010110;
				18'b001101111000001011: oled_data = 16'b1111011000111010;
				18'b001101111010001011: oled_data = 16'b1001010000010000;
				18'b001101111100001011: oled_data = 16'b0100101000000110;
				18'b001101111110001011: oled_data = 16'b0100101001000111;
				18'b001110000000001011: oled_data = 16'b0101101011001001;
				18'b001110000010001011: oled_data = 16'b0110001100001010;
				18'b001110000100001011: oled_data = 16'b0101101011101010;
				18'b001110000110001011: oled_data = 16'b0010100101100101;
				18'b001110001000001011: oled_data = 16'b0001100011100011;
				18'b001110001010001011: oled_data = 16'b0010000100100100;
				18'b001110001100001011: oled_data = 16'b0010000101000101;
				18'b001110001110001011: oled_data = 16'b0010000101000101;
				18'b001110010000001011: oled_data = 16'b0010000101100110;
				18'b001110010010001011: oled_data = 16'b0011000110000110;
				18'b001110010100001011: oled_data = 16'b0011100111000110;
				18'b001110010110001011: oled_data = 16'b0100001000000110;
				18'b001110011000001011: oled_data = 16'b0101001000100111;
				18'b001110011010001011: oled_data = 16'b0101101001100111;
				18'b001110011100001011: oled_data = 16'b0111001011001000;
				18'b001110011110001011: oled_data = 16'b1010001110001100;
				18'b001110100000001011: oled_data = 16'b1100010001010000;
				18'b001110100010001011: oled_data = 16'b1101110010110010;
				18'b001110100100001011: oled_data = 16'b1101110001010001;
				18'b001110100110001011: oled_data = 16'b1100101101101110;
				18'b001100011000001100: oled_data = 16'b0110001010101000;
				18'b001100011010001100: oled_data = 16'b0110001010001000;
				18'b001100011100001100: oled_data = 16'b1010010001010001;
				18'b001100011110001100: oled_data = 16'b1101010010110101;
				18'b001100100000001100: oled_data = 16'b1101010010110101;
				18'b001100100010001100: oled_data = 16'b1101110011010110;
				18'b001100100100001100: oled_data = 16'b1101110011010110;
				18'b001100100110001100: oled_data = 16'b1101010010010100;
				18'b001100101000001100: oled_data = 16'b1101110010110101;
				18'b001100101010001100: oled_data = 16'b1101110011010101;
				18'b001100101100001100: oled_data = 16'b1101110011010101;
				18'b001100101110001100: oled_data = 16'b1101110011010101;
				18'b001100110000001100: oled_data = 16'b1101110011010101;
				18'b001100110010001100: oled_data = 16'b1101110011010101;
				18'b001100110100001100: oled_data = 16'b1101110011010101;
				18'b001100110110001100: oled_data = 16'b1101110011010101;
				18'b001100111000001100: oled_data = 16'b1101110011010110;
				18'b001100111010001100: oled_data = 16'b1101110011010110;
				18'b001100111100001100: oled_data = 16'b1101110011010101;
				18'b001100111110001100: oled_data = 16'b1101110011010101;
				18'b001101000000001100: oled_data = 16'b1101010010010100;
				18'b001101000010001100: oled_data = 16'b1101110011010101;
				18'b001101000100001100: oled_data = 16'b1101110011010101;
				18'b001101000110001100: oled_data = 16'b1101110011010101;
				18'b001101001000001100: oled_data = 16'b1101110011010101;
				18'b001101001010001100: oled_data = 16'b1101110011010101;
				18'b001101001100001100: oled_data = 16'b1101110011010110;
				18'b001101001110001100: oled_data = 16'b1101110011010101;
				18'b001101010000001100: oled_data = 16'b1101110011010101;
				18'b001101010010001100: oled_data = 16'b1101110011010101;
				18'b001101010100001100: oled_data = 16'b1101110011010101;
				18'b001101010110001100: oled_data = 16'b1101110011010101;
				18'b001101011000001100: oled_data = 16'b1101110011010101;
				18'b001101011010001100: oled_data = 16'b1101110011010101;
				18'b001101011100001100: oled_data = 16'b1101110011010101;
				18'b001101011110001100: oled_data = 16'b1101110011010101;
				18'b001101100000001100: oled_data = 16'b1101110011010101;
				18'b001101100010001100: oled_data = 16'b1101110011010101;
				18'b001101100100001100: oled_data = 16'b1101110011010101;
				18'b001101100110001100: oled_data = 16'b1101110011010110;
				18'b001101101000001100: oled_data = 16'b1110010011010110;
				18'b001101101010001100: oled_data = 16'b1101110011010110;
				18'b001101101100001100: oled_data = 16'b1101110011010110;
				18'b001101101110001100: oled_data = 16'b1101110011010101;
				18'b001101110000001100: oled_data = 16'b1101110011010101;
				18'b001101110010001100: oled_data = 16'b1101110011010101;
				18'b001101110100001100: oled_data = 16'b1101110011010101;
				18'b001101110110001100: oled_data = 16'b1101110011010101;
				18'b001101111000001100: oled_data = 16'b1110010100110111;
				18'b001101111010001100: oled_data = 16'b1110011000011001;
				18'b001101111100001100: oled_data = 16'b0111101100101011;
				18'b001101111110001100: oled_data = 16'b0110101100001010;
				18'b001110000000001100: oled_data = 16'b0111101110001011;
				18'b001110000010001100: oled_data = 16'b1000001111101100;
				18'b001110000100001100: oled_data = 16'b0110101101101011;
				18'b001110000110001100: oled_data = 16'b0010000101000100;
				18'b001110001000001100: oled_data = 16'b0001000011000011;
				18'b001110001010001100: oled_data = 16'b0001100100000100;
				18'b001110001100001100: oled_data = 16'b0010000100100101;
				18'b001110001110001100: oled_data = 16'b0010000101000101;
				18'b001110010000001100: oled_data = 16'b0010000101100110;
				18'b001110010010001100: oled_data = 16'b0010100101100110;
				18'b001110010100001100: oled_data = 16'b0010100110000110;
				18'b001110010110001100: oled_data = 16'b0010100110000111;
				18'b001110011000001100: oled_data = 16'b0010100110100111;
				18'b001110011010001100: oled_data = 16'b0110101010101010;
				18'b001110011100001100: oled_data = 16'b1011110001010001;
				18'b001110011110001100: oled_data = 16'b1110010011010100;
				18'b001110100000001100: oled_data = 16'b1101110000110001;
				18'b001110100010001100: oled_data = 16'b1100001100001100;
				18'b001110100100001100: oled_data = 16'b1010101001001001;
				18'b001110100110001100: oled_data = 16'b1010101000001000;
				18'b001100011000001101: oled_data = 16'b1000110010110000;
				18'b001100011010001101: oled_data = 16'b1001010010110001;
				18'b001100011100001101: oled_data = 16'b1100010011110100;
				18'b001100011110001101: oled_data = 16'b1101010001110100;
				18'b001100100000001101: oled_data = 16'b1101110011010110;
				18'b001100100010001101: oled_data = 16'b1101110011010110;
				18'b001100100100001101: oled_data = 16'b1101110011010101;
				18'b001100100110001101: oled_data = 16'b1101010010010100;
				18'b001100101000001101: oled_data = 16'b1101110011010110;
				18'b001100101010001101: oled_data = 16'b1101110011010101;
				18'b001100101100001101: oled_data = 16'b1101110011010101;
				18'b001100101110001101: oled_data = 16'b1101110011010101;
				18'b001100110000001101: oled_data = 16'b1101010010010101;
				18'b001100110010001101: oled_data = 16'b1101110011010110;
				18'b001100110100001101: oled_data = 16'b1101110011010101;
				18'b001100110110001101: oled_data = 16'b1101110011010101;
				18'b001100111000001101: oled_data = 16'b1110010011010110;
				18'b001100111010001101: oled_data = 16'b1110010011010110;
				18'b001100111100001101: oled_data = 16'b1110010011010110;
				18'b001100111110001101: oled_data = 16'b1110010011010110;
				18'b001101000000001101: oled_data = 16'b1101010010010100;
				18'b001101000010001101: oled_data = 16'b1101110010110101;
				18'b001101000100001101: oled_data = 16'b1101110011010101;
				18'b001101000110001101: oled_data = 16'b1101110011010101;
				18'b001101001000001101: oled_data = 16'b1101110011010101;
				18'b001101001010001101: oled_data = 16'b1101110011010101;
				18'b001101001100001101: oled_data = 16'b1110010011010110;
				18'b001101001110001101: oled_data = 16'b1101110011010101;
				18'b001101010000001101: oled_data = 16'b1101110011010101;
				18'b001101010010001101: oled_data = 16'b1101110011010101;
				18'b001101010100001101: oled_data = 16'b1101110011010101;
				18'b001101010110001101: oled_data = 16'b1101110011010101;
				18'b001101011000001101: oled_data = 16'b1101110011010101;
				18'b001101011010001101: oled_data = 16'b1101110011010101;
				18'b001101011100001101: oled_data = 16'b1101110011010101;
				18'b001101011110001101: oled_data = 16'b1101110011010101;
				18'b001101100000001101: oled_data = 16'b1101110011010101;
				18'b001101100010001101: oled_data = 16'b1101110011010101;
				18'b001101100100001101: oled_data = 16'b1101110011010101;
				18'b001101100110001101: oled_data = 16'b1101110011010101;
				18'b001101101000001101: oled_data = 16'b1101110011010101;
				18'b001101101010001101: oled_data = 16'b1101110011010101;
				18'b001101101100001101: oled_data = 16'b1101110011010101;
				18'b001101101110001101: oled_data = 16'b1101110011010101;
				18'b001101110000001101: oled_data = 16'b1101110011010101;
				18'b001101110010001101: oled_data = 16'b1101110011010101;
				18'b001101110100001101: oled_data = 16'b1101110011010101;
				18'b001101110110001101: oled_data = 16'b1101110011010101;
				18'b001101111000001101: oled_data = 16'b1101110011010101;
				18'b001101111010001101: oled_data = 16'b1110110111011001;
				18'b001101111100001101: oled_data = 16'b1011010011110011;
				18'b001101111110001101: oled_data = 16'b0110101011101001;
				18'b001110000000001101: oled_data = 16'b0110101101001010;
				18'b001110000010001101: oled_data = 16'b0110101100101001;
				18'b001110000100001101: oled_data = 16'b0100101001100111;
				18'b001110000110001101: oled_data = 16'b0001100011100011;
				18'b001110001000001101: oled_data = 16'b0001000011000011;
				18'b001110001010001101: oled_data = 16'b0001100011100100;
				18'b001110001100001101: oled_data = 16'b0010000100000100;
				18'b001110001110001101: oled_data = 16'b0010000100100101;
				18'b001110010000001101: oled_data = 16'b0010000101000110;
				18'b001110010010001101: oled_data = 16'b0010000101100110;
				18'b001110010100001101: oled_data = 16'b0010000101100110;
				18'b001110010110001101: oled_data = 16'b0100001000001000;
				18'b001110011000001101: oled_data = 16'b1010101111110000;
				18'b001110011010001101: oled_data = 16'b1110010100010100;
				18'b001110011100001101: oled_data = 16'b1110010010010010;
				18'b001110011110001101: oled_data = 16'b1100001100101101;
				18'b001110100000001101: oled_data = 16'b1011001001001001;
				18'b001110100010001101: oled_data = 16'b1011001000101000;
				18'b001110100100001101: oled_data = 16'b1010101000101000;
				18'b001110100110001101: oled_data = 16'b1010101000001000;
				18'b001100011000001110: oled_data = 16'b0111111000111011;
				18'b001100011010001110: oled_data = 16'b1000110111111000;
				18'b001100011100001110: oled_data = 16'b1100110010010100;
				18'b001100011110001110: oled_data = 16'b1101110010010101;
				18'b001100100000001110: oled_data = 16'b1101110011010110;
				18'b001100100010001110: oled_data = 16'b1101110011010110;
				18'b001100100100001110: oled_data = 16'b1101110010110101;
				18'b001100100110001110: oled_data = 16'b1101010010010100;
				18'b001100101000001110: oled_data = 16'b1101110011010110;
				18'b001100101010001110: oled_data = 16'b1101110011010101;
				18'b001100101100001110: oled_data = 16'b1101110011010110;
				18'b001100101110001110: oled_data = 16'b1101110010010101;
				18'b001100110000001110: oled_data = 16'b1101010010010101;
				18'b001100110010001110: oled_data = 16'b1101110011010110;
				18'b001100110100001110: oled_data = 16'b1101110011010101;
				18'b001100110110001110: oled_data = 16'b1101110011010101;
				18'b001100111000001110: oled_data = 16'b1110010011010110;
				18'b001100111010001110: oled_data = 16'b1110010011010110;
				18'b001100111100001110: oled_data = 16'b1101110011010110;
				18'b001100111110001110: oled_data = 16'b1101110011010110;
				18'b001101000000001110: oled_data = 16'b1101110010110101;
				18'b001101000010001110: oled_data = 16'b1101010001110100;
				18'b001101000100001110: oled_data = 16'b1101110011010110;
				18'b001101000110001110: oled_data = 16'b1101110011010101;
				18'b001101001000001110: oled_data = 16'b1101110011010101;
				18'b001101001010001110: oled_data = 16'b1101110011010101;
				18'b001101001100001110: oled_data = 16'b1101110011010110;
				18'b001101001110001110: oled_data = 16'b1101110011010101;
				18'b001101010000001110: oled_data = 16'b1101110011010101;
				18'b001101010010001110: oled_data = 16'b1101110011010101;
				18'b001101010100001110: oled_data = 16'b1101110011010101;
				18'b001101010110001110: oled_data = 16'b1101110011010101;
				18'b001101011000001110: oled_data = 16'b1101110011010101;
				18'b001101011010001110: oled_data = 16'b1101110011010101;
				18'b001101011100001110: oled_data = 16'b1101110011010101;
				18'b001101011110001110: oled_data = 16'b1101110011010101;
				18'b001101100000001110: oled_data = 16'b1101110011010101;
				18'b001101100010001110: oled_data = 16'b1101110011010101;
				18'b001101100100001110: oled_data = 16'b1101110011010101;
				18'b001101100110001110: oled_data = 16'b1101110011010101;
				18'b001101101000001110: oled_data = 16'b1101110011010101;
				18'b001101101010001110: oled_data = 16'b1101110011010101;
				18'b001101101100001110: oled_data = 16'b1101110011010101;
				18'b001101101110001110: oled_data = 16'b1101110011010101;
				18'b001101110000001110: oled_data = 16'b1101110011010101;
				18'b001101110010001110: oled_data = 16'b1101110011010101;
				18'b001101110100001110: oled_data = 16'b1101110011010101;
				18'b001101110110001110: oled_data = 16'b1101110011010101;
				18'b001101111000001110: oled_data = 16'b1101110011010101;
				18'b001101111010001110: oled_data = 16'b1110010100010110;
				18'b001101111100001110: oled_data = 16'b1110010111111000;
				18'b001101111110001110: oled_data = 16'b0110001011001001;
				18'b001110000000001110: oled_data = 16'b0011100111100110;
				18'b001110000010001110: oled_data = 16'b0011000110100101;
				18'b001110000100001110: oled_data = 16'b0010100101000100;
				18'b001110000110001110: oled_data = 16'b0010000100000100;
				18'b001110001000001110: oled_data = 16'b0001100011100100;
				18'b001110001010001110: oled_data = 16'b0001100011100100;
				18'b001110001100001110: oled_data = 16'b0001100100000100;
				18'b001110001110001110: oled_data = 16'b0010000100100101;
				18'b001110010000001110: oled_data = 16'b0010000101000101;
				18'b001110010010001110: oled_data = 16'b0010000101000101;
				18'b001110010100001110: oled_data = 16'b0110001010001010;
				18'b001110010110001110: oled_data = 16'b1101010010010010;
				18'b001110011000001110: oled_data = 16'b1110110011110100;
				18'b001110011010001110: oled_data = 16'b1101001111001111;
				18'b001110011100001110: oled_data = 16'b1011101010001010;
				18'b001110011110001110: oled_data = 16'b1011001000001000;
				18'b001110100000001110: oled_data = 16'b1011001000101001;
				18'b001110100010001110: oled_data = 16'b1011001000101000;
				18'b001110100100001110: oled_data = 16'b1010101000101000;
				18'b001110100110001110: oled_data = 16'b1010101000001000;
				18'b001100011000001111: oled_data = 16'b1010011011111100;
				18'b001100011010001111: oled_data = 16'b1011010110111000;
				18'b001100011100001111: oled_data = 16'b1101010001110100;
				18'b001100011110001111: oled_data = 16'b1101110011010101;
				18'b001100100000001111: oled_data = 16'b1101110011010101;
				18'b001100100010001111: oled_data = 16'b1101110011010110;
				18'b001100100100001111: oled_data = 16'b1101010001110100;
				18'b001100100110001111: oled_data = 16'b1101110010110101;
				18'b001100101000001111: oled_data = 16'b1101110011010101;
				18'b001100101010001111: oled_data = 16'b1101110011010101;
				18'b001100101100001111: oled_data = 16'b1101110011010110;
				18'b001100101110001111: oled_data = 16'b1101010001010100;
				18'b001100110000001111: oled_data = 16'b1101110010110101;
				18'b001100110010001111: oled_data = 16'b1101110011010101;
				18'b001100110100001111: oled_data = 16'b1101110011010101;
				18'b001100110110001111: oled_data = 16'b1101110011010101;
				18'b001100111000001111: oled_data = 16'b1110010011010110;
				18'b001100111010001111: oled_data = 16'b1110010011010110;
				18'b001100111100001111: oled_data = 16'b1101110011010101;
				18'b001100111110001111: oled_data = 16'b1101110011010101;
				18'b001101000000001111: oled_data = 16'b1101110011010110;
				18'b001101000010001111: oled_data = 16'b1101010001110100;
				18'b001101000100001111: oled_data = 16'b1101110010110101;
				18'b001101000110001111: oled_data = 16'b1101110011010110;
				18'b001101001000001111: oled_data = 16'b1101110011010101;
				18'b001101001010001111: oled_data = 16'b1101110011010101;
				18'b001101001100001111: oled_data = 16'b1101110011010101;
				18'b001101001110001111: oled_data = 16'b1101110011010101;
				18'b001101010000001111: oled_data = 16'b1101110011010101;
				18'b001101010010001111: oled_data = 16'b1101110011010101;
				18'b001101010100001111: oled_data = 16'b1101110011010101;
				18'b001101010110001111: oled_data = 16'b1101110011010101;
				18'b001101011000001111: oled_data = 16'b1101110011010101;
				18'b001101011010001111: oled_data = 16'b1101110011010101;
				18'b001101011100001111: oled_data = 16'b1101110011010101;
				18'b001101011110001111: oled_data = 16'b1110010011110110;
				18'b001101100000001111: oled_data = 16'b1110010011110110;
				18'b001101100010001111: oled_data = 16'b1101110011010101;
				18'b001101100100001111: oled_data = 16'b1101110011010101;
				18'b001101100110001111: oled_data = 16'b1101110011010101;
				18'b001101101000001111: oled_data = 16'b1101110011010101;
				18'b001101101010001111: oled_data = 16'b1101110011010101;
				18'b001101101100001111: oled_data = 16'b1101110011010101;
				18'b001101101110001111: oled_data = 16'b1101110011010101;
				18'b001101110000001111: oled_data = 16'b1101110011010101;
				18'b001101110010001111: oled_data = 16'b1101110011010101;
				18'b001101110100001111: oled_data = 16'b1101110011010101;
				18'b001101110110001111: oled_data = 16'b1101110011010101;
				18'b001101111000001111: oled_data = 16'b1101110011010110;
				18'b001101111010001111: oled_data = 16'b1101110011010101;
				18'b001101111100001111: oled_data = 16'b1110010110010111;
				18'b001101111110001111: oled_data = 16'b1010010001110001;
				18'b001110000000001111: oled_data = 16'b0010000100000100;
				18'b001110000010001111: oled_data = 16'b0010000101000101;
				18'b001110000100001111: oled_data = 16'b0010000100100101;
				18'b001110000110001111: oled_data = 16'b0010000100100100;
				18'b001110001000001111: oled_data = 16'b0001100011100100;
				18'b001110001010001111: oled_data = 16'b0001100011100100;
				18'b001110001100001111: oled_data = 16'b0001100100000100;
				18'b001110001110001111: oled_data = 16'b0001100100100101;
				18'b001110010000001111: oled_data = 16'b0001100100100101;
				18'b001110010010001111: oled_data = 16'b0111101100001100;
				18'b001110010100001111: oled_data = 16'b1110010100010100;
				18'b001110010110001111: oled_data = 16'b1110010010110010;
				18'b001110011000001111: oled_data = 16'b1100001100001100;
				18'b001110011010001111: oled_data = 16'b1011001000101001;
				18'b001110011100001111: oled_data = 16'b1011001000101001;
				18'b001110011110001111: oled_data = 16'b1011001000101001;
				18'b001110100000001111: oled_data = 16'b1011001000101001;
				18'b001110100010001111: oled_data = 16'b1011001000101000;
				18'b001110100100001111: oled_data = 16'b1010101000101000;
				18'b001110100110001111: oled_data = 16'b1010101000001000;
				18'b001100011000010000: oled_data = 16'b1011011011111100;
				18'b001100011010010000: oled_data = 16'b1100010100010110;
				18'b001100011100010000: oled_data = 16'b1101110010010101;
				18'b001100011110010000: oled_data = 16'b1101110011010110;
				18'b001100100000010000: oled_data = 16'b1101110011010101;
				18'b001100100010010000: oled_data = 16'b1101110011010101;
				18'b001100100100010000: oled_data = 16'b1101010001110100;
				18'b001100100110010000: oled_data = 16'b1101110011010101;
				18'b001100101000010000: oled_data = 16'b1101110011010101;
				18'b001100101010010000: oled_data = 16'b1101110011010101;
				18'b001100101100010000: oled_data = 16'b1101110010110101;
				18'b001100101110010000: oled_data = 16'b1100110000010011;
				18'b001100110000010000: oled_data = 16'b1110010011010110;
				18'b001100110010010000: oled_data = 16'b1101110011010101;
				18'b001100110100010000: oled_data = 16'b1101110011010101;
				18'b001100110110010000: oled_data = 16'b1101110011010101;
				18'b001100111000010000: oled_data = 16'b1110010011010110;
				18'b001100111010010000: oled_data = 16'b1110010011010110;
				18'b001100111100010000: oled_data = 16'b1101110011010101;
				18'b001100111110010000: oled_data = 16'b1101110011010101;
				18'b001101000000010000: oled_data = 16'b1101110011010101;
				18'b001101000010010000: oled_data = 16'b1101110010110101;
				18'b001101000100010000: oled_data = 16'b1101010010010100;
				18'b001101000110010000: oled_data = 16'b1110010011010110;
				18'b001101001000010000: oled_data = 16'b1101110011010101;
				18'b001101001010010000: oled_data = 16'b1101110011010101;
				18'b001101001100010000: oled_data = 16'b1101110011010101;
				18'b001101001110010000: oled_data = 16'b1101110011010101;
				18'b001101010000010000: oled_data = 16'b1101110011010101;
				18'b001101010010010000: oled_data = 16'b1101110011010101;
				18'b001101010100010000: oled_data = 16'b1101110011010101;
				18'b001101010110010000: oled_data = 16'b1101110011010101;
				18'b001101011000010000: oled_data = 16'b1101110011010101;
				18'b001101011010010000: oled_data = 16'b1101110011010101;
				18'b001101011100010000: oled_data = 16'b1101110011010101;
				18'b001101011110010000: oled_data = 16'b1101110011010110;
				18'b001101100000010000: oled_data = 16'b1110010011110110;
				18'b001101100010010000: oled_data = 16'b1101110011010101;
				18'b001101100100010000: oled_data = 16'b1101110011010101;
				18'b001101100110010000: oled_data = 16'b1101110011010101;
				18'b001101101000010000: oled_data = 16'b1101110011010101;
				18'b001101101010010000: oled_data = 16'b1101110011010101;
				18'b001101101100010000: oled_data = 16'b1101110011010101;
				18'b001101101110010000: oled_data = 16'b1101110011010101;
				18'b001101110000010000: oled_data = 16'b1101110011010101;
				18'b001101110010010000: oled_data = 16'b1101110011010101;
				18'b001101110100010000: oled_data = 16'b1101110011010101;
				18'b001101110110010000: oled_data = 16'b1101110011010101;
				18'b001101111000010000: oled_data = 16'b1101110011010110;
				18'b001101111010010000: oled_data = 16'b1101110011010110;
				18'b001101111100010000: oled_data = 16'b1101110011110110;
				18'b001101111110010000: oled_data = 16'b1110010110010111;
				18'b001110000000010000: oled_data = 16'b0100100111101000;
				18'b001110000010010000: oled_data = 16'b0010000100100100;
				18'b001110000100010000: oled_data = 16'b0011000101100101;
				18'b001110000110010000: oled_data = 16'b0011000101100101;
				18'b001110001000010000: oled_data = 16'b0010000100000100;
				18'b001110001010010000: oled_data = 16'b0001100011100011;
				18'b001110001100010000: oled_data = 16'b0001100100000100;
				18'b001110001110010000: oled_data = 16'b0001100100100101;
				18'b001110010000010000: oled_data = 16'b1000001100101101;
				18'b001110010010010000: oled_data = 16'b1110110100010101;
				18'b001110010100010000: oled_data = 16'b1101110001010001;
				18'b001110010110010000: oled_data = 16'b1011101010101010;
				18'b001110011000010000: oled_data = 16'b1011001000101001;
				18'b001110011010010000: oled_data = 16'b1011001000101001;
				18'b001110011100010000: oled_data = 16'b1011001000101001;
				18'b001110011110010000: oled_data = 16'b1011001000101001;
				18'b001110100000010000: oled_data = 16'b1011001000101001;
				18'b001110100010010000: oled_data = 16'b1011001000101000;
				18'b001110100100010000: oled_data = 16'b1010101000101000;
				18'b001110100110010000: oled_data = 16'b1010101000001000;
				18'b001100011000010001: oled_data = 16'b1000110100110111;
				18'b001100011010010001: oled_data = 16'b1100110010010100;
				18'b001100011100010001: oled_data = 16'b1101110010110101;
				18'b001100011110010001: oled_data = 16'b1101110011010101;
				18'b001100100000010001: oled_data = 16'b1101110011010101;
				18'b001100100010010001: oled_data = 16'b1101110010110101;
				18'b001100100100010001: oled_data = 16'b1101010010010100;
				18'b001100100110010001: oled_data = 16'b1101110011010110;
				18'b001100101000010001: oled_data = 16'b1110010011010110;
				18'b001100101010010001: oled_data = 16'b1101110011010110;
				18'b001100101100010001: oled_data = 16'b1101010010010100;
				18'b001100101110010001: oled_data = 16'b1101010001010100;
				18'b001100110000010001: oled_data = 16'b1110010011010110;
				18'b001100110010010001: oled_data = 16'b1101110011010101;
				18'b001100110100010001: oled_data = 16'b1101110011010101;
				18'b001100110110010001: oled_data = 16'b1101110011010101;
				18'b001100111000010001: oled_data = 16'b1110010011010110;
				18'b001100111010010001: oled_data = 16'b1101110011010110;
				18'b001100111100010001: oled_data = 16'b1101110011010101;
				18'b001100111110010001: oled_data = 16'b1101110011010101;
				18'b001101000000010001: oled_data = 16'b1101110011010101;
				18'b001101000010010001: oled_data = 16'b1101110011010110;
				18'b001101000100010001: oled_data = 16'b1101010010010100;
				18'b001101000110010001: oled_data = 16'b1101110010110101;
				18'b001101001000010001: oled_data = 16'b1101110011010101;
				18'b001101001010010001: oled_data = 16'b1101110011010101;
				18'b001101001100010001: oled_data = 16'b1101110011010110;
				18'b001101001110010001: oled_data = 16'b1101110011010101;
				18'b001101010000010001: oled_data = 16'b1101110011010101;
				18'b001101010010010001: oled_data = 16'b1101110011010101;
				18'b001101010100010001: oled_data = 16'b1101110011010101;
				18'b001101010110010001: oled_data = 16'b1110010011010110;
				18'b001101011000010001: oled_data = 16'b1110010011110110;
				18'b001101011010010001: oled_data = 16'b1101110011010101;
				18'b001101011100010001: oled_data = 16'b1101110011010101;
				18'b001101011110010001: oled_data = 16'b1101110011010101;
				18'b001101100000010001: oled_data = 16'b1101110011010101;
				18'b001101100010010001: oled_data = 16'b1101110011010101;
				18'b001101100100010001: oled_data = 16'b1101110011010101;
				18'b001101100110010001: oled_data = 16'b1101110011010101;
				18'b001101101000010001: oled_data = 16'b1101110011010101;
				18'b001101101010010001: oled_data = 16'b1101110011010101;
				18'b001101101100010001: oled_data = 16'b1101110011010101;
				18'b001101101110010001: oled_data = 16'b1101110011010101;
				18'b001101110000010001: oled_data = 16'b1101110011010101;
				18'b001101110010010001: oled_data = 16'b1101110011010101;
				18'b001101110100010001: oled_data = 16'b1101110011010101;
				18'b001101110110010001: oled_data = 16'b1101110011010101;
				18'b001101111000010001: oled_data = 16'b1101110011010101;
				18'b001101111010010001: oled_data = 16'b1101110011010101;
				18'b001101111100010001: oled_data = 16'b1101110011010101;
				18'b001101111110010001: oled_data = 16'b1110110101010111;
				18'b001110000000010001: oled_data = 16'b1010010000110001;
				18'b001110000010010001: oled_data = 16'b0010100101000101;
				18'b001110000100010001: oled_data = 16'b0011000110000110;
				18'b001110000110010001: oled_data = 16'b0011000110000110;
				18'b001110001000010001: oled_data = 16'b0010100101000101;
				18'b001110001010010001: oled_data = 16'b0001100100000100;
				18'b001110001100010001: oled_data = 16'b0001100100000101;
				18'b001110001110010001: oled_data = 16'b1000101100101101;
				18'b001110010000010001: oled_data = 16'b1110110100110101;
				18'b001110010010010001: oled_data = 16'b1101010000010000;
				18'b001110010100010001: oled_data = 16'b1011001001101010;
				18'b001110010110010001: oled_data = 16'b1011001000101001;
				18'b001110011000010001: oled_data = 16'b1011001001001001;
				18'b001110011010010001: oled_data = 16'b1011001000101001;
				18'b001110011100010001: oled_data = 16'b1011001001001001;
				18'b001110011110010001: oled_data = 16'b1011001000101001;
				18'b001110100000010001: oled_data = 16'b1011001000101001;
				18'b001110100010010001: oled_data = 16'b1011001000101000;
				18'b001110100100010001: oled_data = 16'b1011001000001000;
				18'b001110100110010001: oled_data = 16'b1011001000001000;
				18'b001100011000010010: oled_data = 16'b0111010000010100;
				18'b001100011010010010: oled_data = 16'b1101010010010101;
				18'b001100011100010010: oled_data = 16'b1101110011010101;
				18'b001100011110010010: oled_data = 16'b1101110011010101;
				18'b001100100000010010: oled_data = 16'b1101110011010110;
				18'b001100100010010010: oled_data = 16'b1101110010110101;
				18'b001100100100010010: oled_data = 16'b1101010010010101;
				18'b001100100110010010: oled_data = 16'b1101110011010110;
				18'b001100101000010010: oled_data = 16'b1110010100010110;
				18'b001100101010010010: oled_data = 16'b1101110011010110;
				18'b001100101100010010: oled_data = 16'b1100110001010100;
				18'b001100101110010010: oled_data = 16'b1101110010010101;
				18'b001100110000010010: oled_data = 16'b1101110011010110;
				18'b001100110010010010: oled_data = 16'b1101110011010101;
				18'b001100110100010010: oled_data = 16'b1101110011010101;
				18'b001100110110010010: oled_data = 16'b1101110011010101;
				18'b001100111000010010: oled_data = 16'b1101110011010110;
				18'b001100111010010010: oled_data = 16'b1101110011010110;
				18'b001100111100010010: oled_data = 16'b1101110011010101;
				18'b001100111110010010: oled_data = 16'b1101110011010101;
				18'b001101000000010010: oled_data = 16'b1101110011010101;
				18'b001101000010010010: oled_data = 16'b1101110011010101;
				18'b001101000100010010: oled_data = 16'b1101110010110101;
				18'b001101000110010010: oled_data = 16'b1101010010010100;
				18'b001101001000010010: oled_data = 16'b1101110011010110;
				18'b001101001010010010: oled_data = 16'b1101110011010101;
				18'b001101001100010010: oled_data = 16'b1101110011010110;
				18'b001101001110010010: oled_data = 16'b1101110011010101;
				18'b001101010000010010: oled_data = 16'b1101110011010101;
				18'b001101010010010010: oled_data = 16'b1101110011010101;
				18'b001101010100010010: oled_data = 16'b1101110011010101;
				18'b001101010110010010: oled_data = 16'b1110010011110110;
				18'b001101011000010010: oled_data = 16'b1110110100110111;
				18'b001101011010010010: oled_data = 16'b1101110011010101;
				18'b001101011100010010: oled_data = 16'b1101110011010101;
				18'b001101011110010010: oled_data = 16'b1101110011010101;
				18'b001101100000010010: oled_data = 16'b1101110011010101;
				18'b001101100010010010: oled_data = 16'b1101110011010101;
				18'b001101100100010010: oled_data = 16'b1101110011010101;
				18'b001101100110010010: oled_data = 16'b1101110011010101;
				18'b001101101000010010: oled_data = 16'b1101110011010101;
				18'b001101101010010010: oled_data = 16'b1101110011010101;
				18'b001101101100010010: oled_data = 16'b1101110011010101;
				18'b001101101110010010: oled_data = 16'b1101110011010101;
				18'b001101110000010010: oled_data = 16'b1101110011010101;
				18'b001101110010010010: oled_data = 16'b1101110011010110;
				18'b001101110100010010: oled_data = 16'b1101110011010101;
				18'b001101110110010010: oled_data = 16'b1101110011010101;
				18'b001101111000010010: oled_data = 16'b1101110011010101;
				18'b001101111010010010: oled_data = 16'b1101110011010101;
				18'b001101111100010010: oled_data = 16'b1101110011010101;
				18'b001101111110010010: oled_data = 16'b1110010011010101;
				18'b001110000000010010: oled_data = 16'b1101110100110110;
				18'b001110000010010010: oled_data = 16'b0101101000101001;
				18'b001110000100010010: oled_data = 16'b0010100101000101;
				18'b001110000110010010: oled_data = 16'b0011000110000110;
				18'b001110001000010010: oled_data = 16'b0010000101000101;
				18'b001110001010010010: oled_data = 16'b0001100100000100;
				18'b001110001100010010: oled_data = 16'b0111101011101100;
				18'b001110001110010010: oled_data = 16'b1110110100110100;
				18'b001110010000010010: oled_data = 16'b1101110000110000;
				18'b001110010010010010: oled_data = 16'b1011001001101010;
				18'b001110010100010010: oled_data = 16'b1011001001001001;
				18'b001110010110010010: oled_data = 16'b1011001001001001;
				18'b001110011000010010: oled_data = 16'b1011001001001001;
				18'b001110011010010010: oled_data = 16'b1011001000101001;
				18'b001110011100010010: oled_data = 16'b1011001001001001;
				18'b001110011110010010: oled_data = 16'b1011001000101001;
				18'b001110100000010010: oled_data = 16'b1011001000101001;
				18'b001110100010010010: oled_data = 16'b1011001000101000;
				18'b001110100100010010: oled_data = 16'b1011001000101000;
				18'b001110100110010010: oled_data = 16'b1011001000001000;
				18'b001100011000010011: oled_data = 16'b1000110000010100;
				18'b001100011010010011: oled_data = 16'b1101010010110101;
				18'b001100011100010011: oled_data = 16'b1101110011010101;
				18'b001100011110010011: oled_data = 16'b1101110011010110;
				18'b001100100000010011: oled_data = 16'b1101110011010110;
				18'b001100100010010011: oled_data = 16'b1101110010010101;
				18'b001100100100010011: oled_data = 16'b1101010010010101;
				18'b001100100110010011: oled_data = 16'b1101110011110110;
				18'b001100101000010011: oled_data = 16'b1101110100010110;
				18'b001100101010010011: oled_data = 16'b1101110011110101;
				18'b001100101100010011: oled_data = 16'b1100110001010011;
				18'b001100101110010011: oled_data = 16'b1101110010110101;
				18'b001100110000010011: oled_data = 16'b1101110011010110;
				18'b001100110010010011: oled_data = 16'b1101110011010101;
				18'b001100110100010011: oled_data = 16'b1101110011010101;
				18'b001100110110010011: oled_data = 16'b1110010100010110;
				18'b001100111000010011: oled_data = 16'b1110010011110110;
				18'b001100111010010011: oled_data = 16'b1110010011010110;
				18'b001100111100010011: oled_data = 16'b1101110011010101;
				18'b001100111110010011: oled_data = 16'b1101110011010101;
				18'b001101000000010011: oled_data = 16'b1101110011010101;
				18'b001101000010010011: oled_data = 16'b1101110011010101;
				18'b001101000100010011: oled_data = 16'b1101110011010101;
				18'b001101000110010011: oled_data = 16'b1101010001010100;
				18'b001101001000010011: oled_data = 16'b1101110011010101;
				18'b001101001010010011: oled_data = 16'b1101110011010101;
				18'b001101001100010011: oled_data = 16'b1101110011010101;
				18'b001101001110010011: oled_data = 16'b1101110011010101;
				18'b001101010000010011: oled_data = 16'b1101110011010101;
				18'b001101010010010011: oled_data = 16'b1101110010110101;
				18'b001101010100010011: oled_data = 16'b1101110011010101;
				18'b001101010110010011: oled_data = 16'b1101110011010101;
				18'b001101011000010011: oled_data = 16'b1110010011110110;
				18'b001101011010010011: oled_data = 16'b1101110011010110;
				18'b001101011100010011: oled_data = 16'b1101110011010101;
				18'b001101011110010011: oled_data = 16'b1101110011010101;
				18'b001101100000010011: oled_data = 16'b1101110011010101;
				18'b001101100010010011: oled_data = 16'b1101110011010101;
				18'b001101100100010011: oled_data = 16'b1101110011010101;
				18'b001101100110010011: oled_data = 16'b1101110011010101;
				18'b001101101000010011: oled_data = 16'b1101110011010101;
				18'b001101101010010011: oled_data = 16'b1101110011010101;
				18'b001101101100010011: oled_data = 16'b1101110011010101;
				18'b001101101110010011: oled_data = 16'b1101110011010101;
				18'b001101110000010011: oled_data = 16'b1101110011010101;
				18'b001101110010010011: oled_data = 16'b1110010011010110;
				18'b001101110100010011: oled_data = 16'b1101110011010101;
				18'b001101110110010011: oled_data = 16'b1101110011010101;
				18'b001101111000010011: oled_data = 16'b1101110011010101;
				18'b001101111010010011: oled_data = 16'b1101110011010101;
				18'b001101111100010011: oled_data = 16'b1101110011010101;
				18'b001101111110010011: oled_data = 16'b1101110011010101;
				18'b001110000000010011: oled_data = 16'b1110010011110110;
				18'b001110000010010011: oled_data = 16'b1010101111010001;
				18'b001110000100010011: oled_data = 16'b0011000101100101;
				18'b001110000110010011: oled_data = 16'b0011000101100110;
				18'b001110001000010011: oled_data = 16'b0010000100100101;
				18'b001110001010010011: oled_data = 16'b0110101010101011;
				18'b001110001100010011: oled_data = 16'b1110010100010100;
				18'b001110001110010011: oled_data = 16'b1101110001010001;
				18'b001110010000010011: oled_data = 16'b1011001010001010;
				18'b001110010010010011: oled_data = 16'b1011001001001001;
				18'b001110010100010011: oled_data = 16'b1011001001001001;
				18'b001110010110010011: oled_data = 16'b1011001001001001;
				18'b001110011000010011: oled_data = 16'b1011001001001001;
				18'b001110011010010011: oled_data = 16'b1011001000101001;
				18'b001110011100010011: oled_data = 16'b1011001001001001;
				18'b001110011110010011: oled_data = 16'b1011001000101001;
				18'b001110100000010011: oled_data = 16'b1011001000101001;
				18'b001110100010010011: oled_data = 16'b1011001000101001;
				18'b001110100100010011: oled_data = 16'b1011001000101000;
				18'b001110100110010011: oled_data = 16'b1011001000001000;
				18'b001100011000010100: oled_data = 16'b1010110000110100;
				18'b001100011010010100: oled_data = 16'b1101110011010101;
				18'b001100011100010100: oled_data = 16'b1101110010110101;
				18'b001100011110010100: oled_data = 16'b1101110011010101;
				18'b001100100000010100: oled_data = 16'b1110010011010110;
				18'b001100100010010100: oled_data = 16'b1101010001010100;
				18'b001100100100010100: oled_data = 16'b1101010010010100;
				18'b001100100110010100: oled_data = 16'b1110010011110110;
				18'b001100101000010100: oled_data = 16'b1101110011110110;
				18'b001100101010010100: oled_data = 16'b1101010011010101;
				18'b001100101100010100: oled_data = 16'b1100110001110100;
				18'b001100101110010100: oled_data = 16'b1101110010110101;
				18'b001100110000010100: oled_data = 16'b1101110011010101;
				18'b001100110010010100: oled_data = 16'b1101110011010101;
				18'b001100110100010100: oled_data = 16'b1101110011010101;
				18'b001100110110010100: oled_data = 16'b1110110110111000;
				18'b001100111000010100: oled_data = 16'b1110010100010110;
				18'b001100111010010100: oled_data = 16'b1110010011010110;
				18'b001100111100010100: oled_data = 16'b1101110011010101;
				18'b001100111110010100: oled_data = 16'b1101110011010101;
				18'b001101000000010100: oled_data = 16'b1101110011010101;
				18'b001101000010010100: oled_data = 16'b1101110011010101;
				18'b001101000100010100: oled_data = 16'b1101110011010110;
				18'b001101000110010100: oled_data = 16'b1101010001110100;
				18'b001101001000010100: oled_data = 16'b1101010010010100;
				18'b001101001010010100: oled_data = 16'b1101110011010110;
				18'b001101001100010100: oled_data = 16'b1101110011010101;
				18'b001101001110010100: oled_data = 16'b1101110011010101;
				18'b001101010000010100: oled_data = 16'b1101110011010101;
				18'b001101010010010100: oled_data = 16'b1101010010010100;
				18'b001101010100010100: oled_data = 16'b1101110011010101;
				18'b001101010110010100: oled_data = 16'b1101110011010101;
				18'b001101011000010100: oled_data = 16'b1101110011010101;
				18'b001101011010010100: oled_data = 16'b1101110011010101;
				18'b001101011100010100: oled_data = 16'b1101110011010101;
				18'b001101011110010100: oled_data = 16'b1101110011010101;
				18'b001101100000010100: oled_data = 16'b1101110011010110;
				18'b001101100010010100: oled_data = 16'b1101110011010101;
				18'b001101100100010100: oled_data = 16'b1101110011010101;
				18'b001101100110010100: oled_data = 16'b1101110011010101;
				18'b001101101000010100: oled_data = 16'b1101110011010101;
				18'b001101101010010100: oled_data = 16'b1101110011010101;
				18'b001101101100010100: oled_data = 16'b1101110011010101;
				18'b001101101110010100: oled_data = 16'b1101110011010101;
				18'b001101110000010100: oled_data = 16'b1101110011010101;
				18'b001101110010010100: oled_data = 16'b1101110011010101;
				18'b001101110100010100: oled_data = 16'b1101110011010101;
				18'b001101110110010100: oled_data = 16'b1101110011010101;
				18'b001101111000010100: oled_data = 16'b1101110011010101;
				18'b001101111010010100: oled_data = 16'b1101110010110101;
				18'b001101111100010100: oled_data = 16'b1101010010010101;
				18'b001101111110010100: oled_data = 16'b1101110011010110;
				18'b001110000000010100: oled_data = 16'b1110010011010110;
				18'b001110000010010100: oled_data = 16'b1101110100010110;
				18'b001110000100010100: oled_data = 16'b0110101010101011;
				18'b001110000110010100: oled_data = 16'b0010100100100101;
				18'b001110001000010100: oled_data = 16'b0101001000101001;
				18'b001110001010010100: oled_data = 16'b1101010011010100;
				18'b001110001100010100: oled_data = 16'b1110010010110011;
				18'b001110001110010100: oled_data = 16'b1011101010101011;
				18'b001110010000010100: oled_data = 16'b1011001001001001;
				18'b001110010010010100: oled_data = 16'b1011101001001001;
				18'b001110010100010100: oled_data = 16'b1011001001001001;
				18'b001110010110010100: oled_data = 16'b1011001001001001;
				18'b001110011000010100: oled_data = 16'b1011001001001001;
				18'b001110011010010100: oled_data = 16'b1011001000101001;
				18'b001110011100010100: oled_data = 16'b1011001001001001;
				18'b001110011110010100: oled_data = 16'b1011001000101001;
				18'b001110100000010100: oled_data = 16'b1010101000001000;
				18'b001110100010010100: oled_data = 16'b1011001000101001;
				18'b001110100100010100: oled_data = 16'b1011001000101000;
				18'b001110100110010100: oled_data = 16'b1011001000001000;
				18'b001100011000010101: oled_data = 16'b1100010001110101;
				18'b001100011010010101: oled_data = 16'b1101110011010110;
				18'b001100011100010101: oled_data = 16'b1101010010010100;
				18'b001100011110010101: oled_data = 16'b1101110011010110;
				18'b001100100000010101: oled_data = 16'b1101110011010110;
				18'b001100100010010101: oled_data = 16'b1100110000110011;
				18'b001100100100010101: oled_data = 16'b1101010010010101;
				18'b001100100110010101: oled_data = 16'b1110010011010110;
				18'b001100101000010101: oled_data = 16'b1101110011010110;
				18'b001100101010010101: oled_data = 16'b1101010010110100;
				18'b001100101100010101: oled_data = 16'b1100010010010010;
				18'b001100101110010101: oled_data = 16'b1101110010010101;
				18'b001100110000010101: oled_data = 16'b1101110011010101;
				18'b001100110010010101: oled_data = 16'b1101110011010101;
				18'b001100110100010101: oled_data = 16'b1101110011010101;
				18'b001100110110010101: oled_data = 16'b1110010101111000;
				18'b001100111000010101: oled_data = 16'b1110010100010110;
				18'b001100111010010101: oled_data = 16'b1101110011010101;
				18'b001100111100010101: oled_data = 16'b1101110011010101;
				18'b001100111110010101: oled_data = 16'b1101110011010101;
				18'b001101000000010101: oled_data = 16'b1101110011010101;
				18'b001101000010010101: oled_data = 16'b1101110011010101;
				18'b001101000100010101: oled_data = 16'b1101110011010101;
				18'b001101000110010101: oled_data = 16'b1101110010110101;
				18'b001101001000010101: oled_data = 16'b1100110000110011;
				18'b001101001010010101: oled_data = 16'b1101110011010110;
				18'b001101001100010101: oled_data = 16'b1101110011010101;
				18'b001101001110010101: oled_data = 16'b1101110011010101;
				18'b001101010000010101: oled_data = 16'b1101110011010110;
				18'b001101010010010101: oled_data = 16'b1101010010110101;
				18'b001101010100010101: oled_data = 16'b1101010010110101;
				18'b001101010110010101: oled_data = 16'b1101110011010110;
				18'b001101011000010101: oled_data = 16'b1101110011010101;
				18'b001101011010010101: oled_data = 16'b1101110011010101;
				18'b001101011100010101: oled_data = 16'b1101110011010110;
				18'b001101011110010101: oled_data = 16'b1101010010010100;
				18'b001101100000010101: oled_data = 16'b1101110010010101;
				18'b001101100010010101: oled_data = 16'b1101110011010110;
				18'b001101100100010101: oled_data = 16'b1101110011010101;
				18'b001101100110010101: oled_data = 16'b1101110011010101;
				18'b001101101000010101: oled_data = 16'b1101110011010101;
				18'b001101101010010101: oled_data = 16'b1101110011010101;
				18'b001101101100010101: oled_data = 16'b1101110011010101;
				18'b001101101110010101: oled_data = 16'b1101110011010101;
				18'b001101110000010101: oled_data = 16'b1101110011010101;
				18'b001101110010010101: oled_data = 16'b1101110011010101;
				18'b001101110100010101: oled_data = 16'b1101110011010101;
				18'b001101110110010101: oled_data = 16'b1101110011010101;
				18'b001101111000010101: oled_data = 16'b1101110011010101;
				18'b001101111010010101: oled_data = 16'b1101110011010101;
				18'b001101111100010101: oled_data = 16'b1101010010010100;
				18'b001101111110010101: oled_data = 16'b1101010010010100;
				18'b001110000000010101: oled_data = 16'b1101110011010110;
				18'b001110000010010101: oled_data = 16'b1110010011110110;
				18'b001110000100010101: oled_data = 16'b1100110010010100;
				18'b001110000110010101: oled_data = 16'b0110001000001001;
				18'b001110001000010101: oled_data = 16'b1011110001010001;
				18'b001110001010010101: oled_data = 16'b1110110100010100;
				18'b001110001100010101: oled_data = 16'b1100001100101101;
				18'b001110001110010101: oled_data = 16'b1011001000101001;
				18'b001110010000010101: oled_data = 16'b1011101001001001;
				18'b001110010010010101: oled_data = 16'b1011101000101001;
				18'b001110010100010101: oled_data = 16'b1011001001001001;
				18'b001110010110010101: oled_data = 16'b1011001001001001;
				18'b001110011000010101: oled_data = 16'b1011001001001001;
				18'b001110011010010101: oled_data = 16'b1011001001001001;
				18'b001110011100010101: oled_data = 16'b1011001000101001;
				18'b001110011110010101: oled_data = 16'b1010001000001000;
				18'b001110100000010101: oled_data = 16'b1010101000001000;
				18'b001110100010010101: oled_data = 16'b1011001000101001;
				18'b001110100100010101: oled_data = 16'b1011001000101000;
				18'b001110100110010101: oled_data = 16'b1011001000001000;
				18'b001100011000010110: oled_data = 16'b1101010001110101;
				18'b001100011010010110: oled_data = 16'b1101110011010101;
				18'b001100011100010110: oled_data = 16'b1100110000110011;
				18'b001100011110010110: oled_data = 16'b1110010011010110;
				18'b001100100000010110: oled_data = 16'b1110010011010110;
				18'b001100100010010110: oled_data = 16'b1100110000010011;
				18'b001100100100010110: oled_data = 16'b1101010010010101;
				18'b001100100110010110: oled_data = 16'b1101110011010110;
				18'b001100101000010110: oled_data = 16'b1101110011010110;
				18'b001100101010010110: oled_data = 16'b1101010011010101;
				18'b001100101100010110: oled_data = 16'b1100110010110011;
				18'b001100101110010110: oled_data = 16'b1101110010010101;
				18'b001100110000010110: oled_data = 16'b1101110010110101;
				18'b001100110010010110: oled_data = 16'b1101110010110101;
				18'b001100110100010110: oled_data = 16'b1101110011010101;
				18'b001100110110010110: oled_data = 16'b1101110100010110;
				18'b001100111000010110: oled_data = 16'b1101110011110110;
				18'b001100111010010110: oled_data = 16'b1101110011010101;
				18'b001100111100010110: oled_data = 16'b1101110011010101;
				18'b001100111110010110: oled_data = 16'b1101110011010101;
				18'b001101000000010110: oled_data = 16'b1101110011010101;
				18'b001101000010010110: oled_data = 16'b1101110011010101;
				18'b001101000100010110: oled_data = 16'b1101110011010101;
				18'b001101000110010110: oled_data = 16'b1101110011010110;
				18'b001101001000010110: oled_data = 16'b1100110000110011;
				18'b001101001010010110: oled_data = 16'b1101110010110101;
				18'b001101001100010110: oled_data = 16'b1101110011010101;
				18'b001101001110010110: oled_data = 16'b1101110011010101;
				18'b001101010000010110: oled_data = 16'b1101110011010101;
				18'b001101010010010110: oled_data = 16'b1101110011010101;
				18'b001101010100010110: oled_data = 16'b1101010001010100;
				18'b001101010110010110: oled_data = 16'b1101110011010110;
				18'b001101011000010110: oled_data = 16'b1101110011010101;
				18'b001101011010010110: oled_data = 16'b1101110011010101;
				18'b001101011100010110: oled_data = 16'b1101110011010101;
				18'b001101011110010110: oled_data = 16'b1101110011010110;
				18'b001101100000010110: oled_data = 16'b1101110010010101;
				18'b001101100010010110: oled_data = 16'b1101010010010100;
				18'b001101100100010110: oled_data = 16'b1101110010110101;
				18'b001101100110010110: oled_data = 16'b1101110011010101;
				18'b001101101000010110: oled_data = 16'b1101110011010110;
				18'b001101101010010110: oled_data = 16'b1101110011010110;
				18'b001101101100010110: oled_data = 16'b1101110011010101;
				18'b001101101110010110: oled_data = 16'b1101110011010101;
				18'b001101110000010110: oled_data = 16'b1101110011010101;
				18'b001101110010010110: oled_data = 16'b1101110011010101;
				18'b001101110100010110: oled_data = 16'b1101110011010101;
				18'b001101110110010110: oled_data = 16'b1101110011010110;
				18'b001101111000010110: oled_data = 16'b1101110011010101;
				18'b001101111010010110: oled_data = 16'b1101110011010101;
				18'b001101111100010110: oled_data = 16'b1101110011010110;
				18'b001101111110010110: oled_data = 16'b1101010010010100;
				18'b001110000000010110: oled_data = 16'b1101010001110100;
				18'b001110000010010110: oled_data = 16'b1101110011010110;
				18'b001110000100010110: oled_data = 16'b1101110011010101;
				18'b001110000110010110: oled_data = 16'b1101010010010011;
				18'b001110001000010110: oled_data = 16'b1110110100010100;
				18'b001110001010010110: oled_data = 16'b1101001111101111;
				18'b001110001100010110: oled_data = 16'b1011001001001001;
				18'b001110001110010110: oled_data = 16'b1011101001001001;
				18'b001110010000010110: oled_data = 16'b1011101001001001;
				18'b001110010010010110: oled_data = 16'b1011101001001001;
				18'b001110010100010110: oled_data = 16'b1011001001001001;
				18'b001110010110010110: oled_data = 16'b1011001001001001;
				18'b001110011000010110: oled_data = 16'b1011001001001001;
				18'b001110011010010110: oled_data = 16'b1010101000101000;
				18'b001110011100010110: oled_data = 16'b1010001000001000;
				18'b001110011110010110: oled_data = 16'b1011001000101001;
				18'b001110100000010110: oled_data = 16'b1011001000101001;
				18'b001110100010010110: oled_data = 16'b1011001000101001;
				18'b001110100100010110: oled_data = 16'b1011001000101000;
				18'b001110100110010110: oled_data = 16'b1011001000001000;
				18'b001100011000010111: oled_data = 16'b1101110010010101;
				18'b001100011010010111: oled_data = 16'b1101010010110100;
				18'b001100011100010111: oled_data = 16'b1100110001110100;
				18'b001100011110010111: oled_data = 16'b1110010011110110;
				18'b001100100000010111: oled_data = 16'b1101110011010110;
				18'b001100100010010111: oled_data = 16'b1100110000010011;
				18'b001100100100010111: oled_data = 16'b1101110010110101;
				18'b001100100110010111: oled_data = 16'b1101110011010110;
				18'b001100101000010111: oled_data = 16'b1101110011010101;
				18'b001100101010010111: oled_data = 16'b1101110100010101;
				18'b001100101100010111: oled_data = 16'b1101010100010101;
				18'b001100101110010111: oled_data = 16'b1101110010110101;
				18'b001100110000010111: oled_data = 16'b1101110010110101;
				18'b001100110010010111: oled_data = 16'b1101010010010101;
				18'b001100110100010111: oled_data = 16'b1101110011010110;
				18'b001100110110010111: oled_data = 16'b1101110011010101;
				18'b001100111000010111: oled_data = 16'b1101110011010101;
				18'b001100111010010111: oled_data = 16'b1101110011010101;
				18'b001100111100010111: oled_data = 16'b1101110011010101;
				18'b001100111110010111: oled_data = 16'b1101110011010101;
				18'b001101000000010111: oled_data = 16'b1101110011010101;
				18'b001101000010010111: oled_data = 16'b1101010010010101;
				18'b001101000100010111: oled_data = 16'b1101110011010101;
				18'b001101000110010111: oled_data = 16'b1101110011010110;
				18'b001101001000010111: oled_data = 16'b1101010001110100;
				18'b001101001010010111: oled_data = 16'b1100110001010100;
				18'b001101001100010111: oled_data = 16'b1101110011010110;
				18'b001101001110010111: oled_data = 16'b1101110011010101;
				18'b001101010000010111: oled_data = 16'b1110010011010101;
				18'b001101010010010111: oled_data = 16'b1110010011010110;
				18'b001101010100010111: oled_data = 16'b1100110001010011;
				18'b001101010110010111: oled_data = 16'b1101010010110101;
				18'b001101011000010111: oled_data = 16'b1101110011010101;
				18'b001101011010010111: oled_data = 16'b1101110011010101;
				18'b001101011100010111: oled_data = 16'b1110010011010101;
				18'b001101011110010111: oled_data = 16'b1101110011010101;
				18'b001101100000010111: oled_data = 16'b1101110011010110;
				18'b001101100010010111: oled_data = 16'b1101110011010101;
				18'b001101100100010111: oled_data = 16'b1101010010010101;
				18'b001101100110010111: oled_data = 16'b1101010001110100;
				18'b001101101000010111: oled_data = 16'b1101010001110100;
				18'b001101101010010111: oled_data = 16'b1101110010010101;
				18'b001101101100010111: oled_data = 16'b1101110010110101;
				18'b001101101110010111: oled_data = 16'b1101110010110101;
				18'b001101110000010111: oled_data = 16'b1101110010110101;
				18'b001101110010010111: oled_data = 16'b1101110010110101;
				18'b001101110100010111: oled_data = 16'b1101110010010101;
				18'b001101110110010111: oled_data = 16'b1101010001110100;
				18'b001101111000010111: oled_data = 16'b1101110010110101;
				18'b001101111010010111: oled_data = 16'b1101110011010110;
				18'b001101111100010111: oled_data = 16'b1101110011010101;
				18'b001101111110010111: oled_data = 16'b1101110011010110;
				18'b001110000000010111: oled_data = 16'b1101010010010101;
				18'b001110000010010111: oled_data = 16'b1101010001010100;
				18'b001110000100010111: oled_data = 16'b1101010001010011;
				18'b001110000110010111: oled_data = 16'b1110010011110100;
				18'b001110001000010111: oled_data = 16'b1110010010110010;
				18'b001110001010010111: oled_data = 16'b1011101010001010;
				18'b001110001100010111: oled_data = 16'b1011001001001001;
				18'b001110001110010111: oled_data = 16'b1011001001001001;
				18'b001110010000010111: oled_data = 16'b1011001001001001;
				18'b001110010010010111: oled_data = 16'b1011001001001001;
				18'b001110010100010111: oled_data = 16'b1011001001001001;
				18'b001110010110010111: oled_data = 16'b1011001001001001;
				18'b001110011000010111: oled_data = 16'b1011001000101001;
				18'b001110011010010111: oled_data = 16'b1010001000001000;
				18'b001110011100010111: oled_data = 16'b1011001001001001;
				18'b001110011110010111: oled_data = 16'b1011001000101001;
				18'b001110100000010111: oled_data = 16'b1011001000101001;
				18'b001110100010010111: oled_data = 16'b1011001000101001;
				18'b001110100100010111: oled_data = 16'b1011001000101000;
				18'b001110100110010111: oled_data = 16'b1011001000001000;
				18'b001100011000011000: oled_data = 16'b1101110010110101;
				18'b001100011010011000: oled_data = 16'b1101010010010011;
				18'b001100011100011000: oled_data = 16'b1100110010010100;
				18'b001100011110011000: oled_data = 16'b1110010011010110;
				18'b001100100000011000: oled_data = 16'b1101110011010110;
				18'b001100100010011000: oled_data = 16'b1100110000110011;
				18'b001100100100011000: oled_data = 16'b1101110010110101;
				18'b001100100110011000: oled_data = 16'b1101110011010110;
				18'b001100101000011000: oled_data = 16'b1101110010110101;
				18'b001100101010011000: oled_data = 16'b1101010101010110;
				18'b001100101100011000: oled_data = 16'b1101010110010110;
				18'b001100101110011000: oled_data = 16'b1101110010010101;
				18'b001100110000011000: oled_data = 16'b1101110010110101;
				18'b001100110010011000: oled_data = 16'b1101010010010100;
				18'b001100110100011000: oled_data = 16'b1101110011010110;
				18'b001100110110011000: oled_data = 16'b1101110011010101;
				18'b001100111000011000: oled_data = 16'b1101110011010101;
				18'b001100111010011000: oled_data = 16'b1101110011010101;
				18'b001100111100011000: oled_data = 16'b1101110011010101;
				18'b001100111110011000: oled_data = 16'b1101110011010101;
				18'b001101000000011000: oled_data = 16'b1110010011010110;
				18'b001101000010011000: oled_data = 16'b1100110001010011;
				18'b001101000100011000: oled_data = 16'b1101010001110100;
				18'b001101000110011000: oled_data = 16'b1101110011010110;
				18'b001101001000011000: oled_data = 16'b1101110011010101;
				18'b001101001010011000: oled_data = 16'b1100110000110011;
				18'b001101001100011000: oled_data = 16'b1101110011010101;
				18'b001101001110011000: oled_data = 16'b1101110011010101;
				18'b001101010000011000: oled_data = 16'b1110010011010101;
				18'b001101010010011000: oled_data = 16'b1101110011010110;
				18'b001101010100011000: oled_data = 16'b1101010010010100;
				18'b001101010110011000: oled_data = 16'b1100110001010011;
				18'b001101011000011000: oled_data = 16'b1110010011010110;
				18'b001101011010011000: oled_data = 16'b1101110011010101;
				18'b001101011100011000: oled_data = 16'b1110010011010101;
				18'b001101011110011000: oled_data = 16'b1101110011010101;
				18'b001101100000011000: oled_data = 16'b1101110011010101;
				18'b001101100010011000: oled_data = 16'b1101110011010101;
				18'b001101100100011000: oled_data = 16'b1101110011010110;
				18'b001101100110011000: oled_data = 16'b1101110011010110;
				18'b001101101000011000: oled_data = 16'b1101110010110101;
				18'b001101101010011000: oled_data = 16'b1101010010010101;
				18'b001101101100011000: oled_data = 16'b1101010010010100;
				18'b001101101110011000: oled_data = 16'b1101010001110100;
				18'b001101110000011000: oled_data = 16'b1101010001110100;
				18'b001101110010011000: oled_data = 16'b1101010001110100;
				18'b001101110100011000: oled_data = 16'b1101010001010100;
				18'b001101110110011000: oled_data = 16'b1100110000110011;
				18'b001101111000011000: oled_data = 16'b1101110010110101;
				18'b001101111010011000: oled_data = 16'b1101110011010101;
				18'b001101111100011000: oled_data = 16'b1101110011010101;
				18'b001101111110011000: oled_data = 16'b1101110011010101;
				18'b001110000000011000: oled_data = 16'b1101110011010110;
				18'b001110000010011000: oled_data = 16'b1101110010010101;
				18'b001110000100011000: oled_data = 16'b1101010010010010;
				18'b001110000110011000: oled_data = 16'b1110110100010100;
				18'b001110001000011000: oled_data = 16'b1100101101101101;
				18'b001110001010011000: oled_data = 16'b1011001000101001;
				18'b001110001100011000: oled_data = 16'b1011001001001001;
				18'b001110001110011000: oled_data = 16'b1011001001001001;
				18'b001110010000011000: oled_data = 16'b1011001001001001;
				18'b001110010010011000: oled_data = 16'b1011001001001001;
				18'b001110010100011000: oled_data = 16'b1011001001001001;
				18'b001110010110011000: oled_data = 16'b1011001000101001;
				18'b001110011000011000: oled_data = 16'b1010101000001000;
				18'b001110011010011000: oled_data = 16'b1011001000101001;
				18'b001110011100011000: oled_data = 16'b1011001001001001;
				18'b001110011110011000: oled_data = 16'b1011001000101001;
				18'b001110100000011000: oled_data = 16'b1011001000101001;
				18'b001110100010011000: oled_data = 16'b1011001000101001;
				18'b001110100100011000: oled_data = 16'b1011001000101000;
				18'b001110100110011000: oled_data = 16'b1010101000001000;
				18'b001100011000011001: oled_data = 16'b1110010011010110;
				18'b001100011010011001: oled_data = 16'b1100010001010000;
				18'b001100011100011001: oled_data = 16'b1100110010010010;
				18'b001100011110011001: oled_data = 16'b1110010011010110;
				18'b001100100000011001: oled_data = 16'b1101110011010110;
				18'b001100100010011001: oled_data = 16'b1100110000010011;
				18'b001100100100011001: oled_data = 16'b1101110010110101;
				18'b001100100110011001: oled_data = 16'b1101110011010110;
				18'b001100101000011001: oled_data = 16'b1101110011010101;
				18'b001100101010011001: oled_data = 16'b1101010110010111;
				18'b001100101100011001: oled_data = 16'b1101110111110111;
				18'b001100101110011001: oled_data = 16'b1101010010010100;
				18'b001100110000011001: oled_data = 16'b1101110010110101;
				18'b001100110010011001: oled_data = 16'b1101010010010100;
				18'b001100110100011001: oled_data = 16'b1101110011010110;
				18'b001100110110011001: oled_data = 16'b1101110011010101;
				18'b001100111000011001: oled_data = 16'b1101110011010101;
				18'b001100111010011001: oled_data = 16'b1101110011010101;
				18'b001100111100011001: oled_data = 16'b1101110011010101;
				18'b001100111110011001: oled_data = 16'b1101110011010101;
				18'b001101000000011001: oled_data = 16'b1101110011010110;
				18'b001101000010011001: oled_data = 16'b1101110010110101;
				18'b001101000100011001: oled_data = 16'b1100110000110011;
				18'b001101000110011001: oled_data = 16'b1101110011010110;
				18'b001101001000011001: oled_data = 16'b1101110011010110;
				18'b001101001010011001: oled_data = 16'b1101010001110100;
				18'b001101001100011001: oled_data = 16'b1101010010010101;
				18'b001101001110011001: oled_data = 16'b1101110011010110;
				18'b001101010000011001: oled_data = 16'b1101110011010101;
				18'b001101010010011001: oled_data = 16'b1101110011010101;
				18'b001101010100011001: oled_data = 16'b1101110011010110;
				18'b001101010110011001: oled_data = 16'b1100110001110100;
				18'b001101011000011001: oled_data = 16'b1101110010110101;
				18'b001101011010011001: oled_data = 16'b1101110011010101;
				18'b001101011100011001: oled_data = 16'b1101110011010101;
				18'b001101011110011001: oled_data = 16'b1101110011010101;
				18'b001101100000011001: oled_data = 16'b1101110011010101;
				18'b001101100010011001: oled_data = 16'b1101110011010101;
				18'b001101100100011001: oled_data = 16'b1101110011010101;
				18'b001101100110011001: oled_data = 16'b1101110011010101;
				18'b001101101000011001: oled_data = 16'b1101110011010101;
				18'b001101101010011001: oled_data = 16'b1101110011010110;
				18'b001101101100011001: oled_data = 16'b1110010011010110;
				18'b001101101110011001: oled_data = 16'b1101110011110110;
				18'b001101110000011001: oled_data = 16'b1110010011110110;
				18'b001101110010011001: oled_data = 16'b1110010011010110;
				18'b001101110100011001: oled_data = 16'b1101010001110100;
				18'b001101110110011001: oled_data = 16'b1101110010110101;
				18'b001101111000011001: oled_data = 16'b1101110011010101;
				18'b001101111010011001: oled_data = 16'b1101110011010101;
				18'b001101111100011001: oled_data = 16'b1101110011010101;
				18'b001101111110011001: oled_data = 16'b1101110011010101;
				18'b001110000000011001: oled_data = 16'b1101110011010101;
				18'b001110000010011001: oled_data = 16'b1101010001110011;
				18'b001110000100011001: oled_data = 16'b1110010011110100;
				18'b001110000110011001: oled_data = 16'b1101110001110001;
				18'b001110001000011001: oled_data = 16'b1011101001101010;
				18'b001110001010011001: oled_data = 16'b1011001001001001;
				18'b001110001100011001: oled_data = 16'b1011001001001001;
				18'b001110001110011001: oled_data = 16'b1011001001001001;
				18'b001110010000011001: oled_data = 16'b1011001001001001;
				18'b001110010010011001: oled_data = 16'b1011001001001001;
				18'b001110010100011001: oled_data = 16'b1011001000101001;
				18'b001110010110011001: oled_data = 16'b1010101000001000;
				18'b001110011000011001: oled_data = 16'b1011001000101001;
				18'b001110011010011001: oled_data = 16'b1011001001001001;
				18'b001110011100011001: oled_data = 16'b1011001000101001;
				18'b001110011110011001: oled_data = 16'b1011001000101001;
				18'b001110100000011001: oled_data = 16'b1011001000101001;
				18'b001110100010011001: oled_data = 16'b1011001000101000;
				18'b001110100100011001: oled_data = 16'b1011001000101000;
				18'b001110100110011001: oled_data = 16'b1010101000101000;
				18'b001100011000011010: oled_data = 16'b1110010011110110;
				18'b001100011010011010: oled_data = 16'b1011110000101110;
				18'b001100011100011010: oled_data = 16'b1100110010010010;
				18'b001100011110011010: oled_data = 16'b1110010011010110;
				18'b001100100000011010: oled_data = 16'b1110010011010110;
				18'b001100100010011010: oled_data = 16'b1100001111110010;
				18'b001100100100011010: oled_data = 16'b1101010001110100;
				18'b001100100110011010: oled_data = 16'b1101110011010110;
				18'b001100101000011010: oled_data = 16'b1101110010110101;
				18'b001100101010011010: oled_data = 16'b1101110110010111;
				18'b001100101100011010: oled_data = 16'b1110111010011010;
				18'b001100101110011010: oled_data = 16'b1101010010110100;
				18'b001100110000011010: oled_data = 16'b1110010011010110;
				18'b001100110010011010: oled_data = 16'b1101010001110100;
				18'b001100110100011010: oled_data = 16'b1101110011010101;
				18'b001100110110011010: oled_data = 16'b1101110011010101;
				18'b001100111000011010: oled_data = 16'b1101110011010101;
				18'b001100111010011010: oled_data = 16'b1101110011010101;
				18'b001100111100011010: oled_data = 16'b1101110011010101;
				18'b001100111110011010: oled_data = 16'b1101110011010101;
				18'b001101000000011010: oled_data = 16'b1101110011010101;
				18'b001101000010011010: oled_data = 16'b1101110011010101;
				18'b001101000100011010: oled_data = 16'b1100110000110011;
				18'b001101000110011010: oled_data = 16'b1101110010110101;
				18'b001101001000011010: oled_data = 16'b1101110011010110;
				18'b001101001010011010: oled_data = 16'b1101110010110101;
				18'b001101001100011010: oled_data = 16'b1100110001010011;
				18'b001101001110011010: oled_data = 16'b1101110011010101;
				18'b001101010000011010: oled_data = 16'b1101110011010101;
				18'b001101010010011010: oled_data = 16'b1101110011010101;
				18'b001101010100011010: oled_data = 16'b1101110011010110;
				18'b001101010110011010: oled_data = 16'b1101010010010100;
				18'b001101011000011010: oled_data = 16'b1100110001110100;
				18'b001101011010011010: oled_data = 16'b1101110011010101;
				18'b001101011100011010: oled_data = 16'b1101110011010101;
				18'b001101011110011010: oled_data = 16'b1101110011010101;
				18'b001101100000011010: oled_data = 16'b1101110011010101;
				18'b001101100010011010: oled_data = 16'b1101110011010101;
				18'b001101100100011010: oled_data = 16'b1101110011010101;
				18'b001101100110011010: oled_data = 16'b1101110011010101;
				18'b001101101000011010: oled_data = 16'b1101110011010101;
				18'b001101101010011010: oled_data = 16'b1101110011010101;
				18'b001101101100011010: oled_data = 16'b1101110011010101;
				18'b001101101110011010: oled_data = 16'b1101110011010110;
				18'b001101110000011010: oled_data = 16'b1101110010110101;
				18'b001101110010011010: oled_data = 16'b1101010001110100;
				18'b001101110100011010: oled_data = 16'b1101110010110101;
				18'b001101110110011010: oled_data = 16'b1101110011010110;
				18'b001101111000011010: oled_data = 16'b1101110011010101;
				18'b001101111010011010: oled_data = 16'b1101110011010101;
				18'b001101111100011010: oled_data = 16'b1110010011010110;
				18'b001101111110011010: oled_data = 16'b1110010011010110;
				18'b001110000000011010: oled_data = 16'b1101110010110100;
				18'b001110000010011010: oled_data = 16'b1101110010110011;
				18'b001110000100011010: oled_data = 16'b1110110100010100;
				18'b001110000110011010: oled_data = 16'b1100101100101101;
				18'b001110001000011010: oled_data = 16'b1011001001001001;
				18'b001110001010011010: oled_data = 16'b1011001001001001;
				18'b001110001100011010: oled_data = 16'b1011001001001001;
				18'b001110001110011010: oled_data = 16'b1011001001001001;
				18'b001110010000011010: oled_data = 16'b1011001001001001;
				18'b001110010010011010: oled_data = 16'b1011001001001001;
				18'b001110010100011010: oled_data = 16'b1010101000001000;
				18'b001110010110011010: oled_data = 16'b1011001000101001;
				18'b001110011000011010: oled_data = 16'b1011001001001001;
				18'b001110011010011010: oled_data = 16'b1011001001001001;
				18'b001110011100011010: oled_data = 16'b1011001000101001;
				18'b001110011110011010: oled_data = 16'b1011001000101001;
				18'b001110100000011010: oled_data = 16'b1011001000101001;
				18'b001110100010011010: oled_data = 16'b1011001000101000;
				18'b001110100100011010: oled_data = 16'b1011001000101000;
				18'b001110100110011010: oled_data = 16'b1010101000101000;
				18'b001100011000011011: oled_data = 16'b1101110011010110;
				18'b001100011010011011: oled_data = 16'b1011010000101100;
				18'b001100011100011011: oled_data = 16'b1100110010110001;
				18'b001100011110011011: oled_data = 16'b1110010011010110;
				18'b001100100000011011: oled_data = 16'b1110010011010110;
				18'b001100100010011011: oled_data = 16'b1100010000010011;
				18'b001100100100011011: oled_data = 16'b1100110001010100;
				18'b001100100110011011: oled_data = 16'b1110010011010110;
				18'b001100101000011011: oled_data = 16'b1101110010110101;
				18'b001100101010011011: oled_data = 16'b1101010110010111;
				18'b001100101100011011: oled_data = 16'b1110011010111010;
				18'b001100101110011011: oled_data = 16'b1101010101110110;
				18'b001100110000011011: oled_data = 16'b1101110011010101;
				18'b001100110010011011: oled_data = 16'b1101010001110100;
				18'b001100110100011011: oled_data = 16'b1101110010110101;
				18'b001100110110011011: oled_data = 16'b1101110011010101;
				18'b001100111000011011: oled_data = 16'b1101110011010101;
				18'b001100111010011011: oled_data = 16'b1101110011010101;
				18'b001100111100011011: oled_data = 16'b1101110011010101;
				18'b001100111110011011: oled_data = 16'b1101110011010101;
				18'b001101000000011011: oled_data = 16'b1101110011010101;
				18'b001101000010011011: oled_data = 16'b1101110011010110;
				18'b001101000100011011: oled_data = 16'b1101010010010100;
				18'b001101000110011011: oled_data = 16'b1101010010010100;
				18'b001101001000011011: oled_data = 16'b1101110011010101;
				18'b001101001010011011: oled_data = 16'b1101110011010101;
				18'b001101001100011011: oled_data = 16'b1100110001110100;
				18'b001101001110011011: oled_data = 16'b1101010011010101;
				18'b001101010000011011: oled_data = 16'b1101110011010110;
				18'b001101010010011011: oled_data = 16'b1101110011010101;
				18'b001101010100011011: oled_data = 16'b1101110011010101;
				18'b001101010110011011: oled_data = 16'b1101110011010101;
				18'b001101011000011011: oled_data = 16'b1101010100010101;
				18'b001101011010011011: oled_data = 16'b1101010011010100;
				18'b001101011100011011: oled_data = 16'b1101110011010101;
				18'b001101011110011011: oled_data = 16'b1101110011010101;
				18'b001101100000011011: oled_data = 16'b1101110011010101;
				18'b001101100010011011: oled_data = 16'b1101110011010110;
				18'b001101100100011011: oled_data = 16'b1101110011010110;
				18'b001101100110011011: oled_data = 16'b1101110011010110;
				18'b001101101000011011: oled_data = 16'b1101110011010110;
				18'b001101101010011011: oled_data = 16'b1101110011010110;
				18'b001101101100011011: oled_data = 16'b1101110011010101;
				18'b001101101110011011: oled_data = 16'b1101010011010101;
				18'b001101110000011011: oled_data = 16'b1011110100010100;
				18'b001101110010011011: oled_data = 16'b1100110100010101;
				18'b001101110100011011: oled_data = 16'b1101110011010101;
				18'b001101110110011011: oled_data = 16'b1101110011010110;
				18'b001101111000011011: oled_data = 16'b1101110011010101;
				18'b001101111010011011: oled_data = 16'b1101010010110101;
				18'b001101111100011011: oled_data = 16'b1101010001110100;
				18'b001101111110011011: oled_data = 16'b1101110010010101;
				18'b001110000000011011: oled_data = 16'b1100110001010010;
				18'b001110000010011011: oled_data = 16'b1110010011110100;
				18'b001110000100011011: oled_data = 16'b1101110001110001;
				18'b001110000110011011: oled_data = 16'b1011101001101010;
				18'b001110001000011011: oled_data = 16'b1011101001001001;
				18'b001110001010011011: oled_data = 16'b1100001011001100;
				18'b001110001100011011: oled_data = 16'b1011101001101010;
				18'b001110001110011011: oled_data = 16'b1011001001001001;
				18'b001110010000011011: oled_data = 16'b1011001001001001;
				18'b001110010010011011: oled_data = 16'b1011001000101000;
				18'b001110010100011011: oled_data = 16'b1010101000101001;
				18'b001110010110011011: oled_data = 16'b1011001001001001;
				18'b001110011000011011: oled_data = 16'b1011001001001001;
				18'b001110011010011011: oled_data = 16'b1011001000101001;
				18'b001110011100011011: oled_data = 16'b1011001000101001;
				18'b001110011110011011: oled_data = 16'b1011001000101001;
				18'b001110100000011011: oled_data = 16'b1011001000101001;
				18'b001110100010011011: oled_data = 16'b1011001000101000;
				18'b001110100100011011: oled_data = 16'b1011001000101000;
				18'b001110100110011011: oled_data = 16'b1010101000101000;
				18'b001100011000011100: oled_data = 16'b1101110011010110;
				18'b001100011010011100: oled_data = 16'b1011010000101011;
				18'b001100011100011100: oled_data = 16'b1100010010010000;
				18'b001100011110011100: oled_data = 16'b1110010011010110;
				18'b001100100000011100: oled_data = 16'b1101110011010110;
				18'b001100100010011100: oled_data = 16'b1100001111110010;
				18'b001100100100011100: oled_data = 16'b1100110000110011;
				18'b001100100110011100: oled_data = 16'b1110010011010110;
				18'b001100101000011100: oled_data = 16'b1101110010110101;
				18'b001100101010011100: oled_data = 16'b1101110110110111;
				18'b001100101100011100: oled_data = 16'b1101111010111001;
				18'b001100101110011100: oled_data = 16'b1101011000011000;
				18'b001100110000011100: oled_data = 16'b1101010010110101;
				18'b001100110010011100: oled_data = 16'b1101110010010101;
				18'b001100110100011100: oled_data = 16'b1101110010110101;
				18'b001100110110011100: oled_data = 16'b1101110011010101;
				18'b001100111000011100: oled_data = 16'b1101110011010101;
				18'b001100111010011100: oled_data = 16'b1101110011010101;
				18'b001100111100011100: oled_data = 16'b1101110011010101;
				18'b001100111110011100: oled_data = 16'b1101110011010101;
				18'b001101000000011100: oled_data = 16'b1101110011010101;
				18'b001101000010011100: oled_data = 16'b1101110011010101;
				18'b001101000100011100: oled_data = 16'b1101010011110101;
				18'b001101000110011100: oled_data = 16'b1100110010110011;
				18'b001101001000011100: oled_data = 16'b1101010010110100;
				18'b001101001010011100: oled_data = 16'b1110010011010101;
				18'b001101001100011100: oled_data = 16'b1101010010010100;
				18'b001101001110011100: oled_data = 16'b1100110010010100;
				18'b001101010000011100: oled_data = 16'b1101110011010101;
				18'b001101010010011100: oled_data = 16'b1101110011010110;
				18'b001101010100011100: oled_data = 16'b1101110011010101;
				18'b001101010110011100: oled_data = 16'b1101110010110101;
				18'b001101011000011100: oled_data = 16'b1101110110010111;
				18'b001101011010011100: oled_data = 16'b1101010110110111;
				18'b001101011100011100: oled_data = 16'b1101010010110101;
				18'b001101011110011100: oled_data = 16'b1101110011010101;
				18'b001101100000011100: oled_data = 16'b1101110011010101;
				18'b001101100010011100: oled_data = 16'b1101010001010100;
				18'b001101100100011100: oled_data = 16'b1100110000110011;
				18'b001101100110011100: oled_data = 16'b1100110001010011;
				18'b001101101000011100: oled_data = 16'b1100110000110011;
				18'b001101101010011100: oled_data = 16'b1100010000010010;
				18'b001101101100011100: oled_data = 16'b1100110000010010;
				18'b001101101110011100: oled_data = 16'b1101010011110101;
				18'b001101110000011100: oled_data = 16'b1111011011111011;
				18'b001101110010011100: oled_data = 16'b1110111011111011;
				18'b001101110100011100: oled_data = 16'b1101010110010110;
				18'b001101110110011100: oled_data = 16'b1101010010010101;
				18'b001101111000011100: oled_data = 16'b1110010011010110;
				18'b001101111010011100: oled_data = 16'b1101110011010101;
				18'b001101111100011100: oled_data = 16'b1101010001110100;
				18'b001101111110011100: oled_data = 16'b1100110000010011;
				18'b001110000000011100: oled_data = 16'b1101010001110010;
				18'b001110000010011100: oled_data = 16'b1110110100010100;
				18'b001110000100011100: oled_data = 16'b1100101101101101;
				18'b001110000110011100: oled_data = 16'b1011001000101001;
				18'b001110001000011100: oled_data = 16'b1011101010001010;
				18'b001110001010011100: oled_data = 16'b1101001110001110;
				18'b001110001100011100: oled_data = 16'b1011001001001010;
				18'b001110001110011100: oled_data = 16'b1011101001001001;
				18'b001110010000011100: oled_data = 16'b1011001001001001;
				18'b001110010010011100: oled_data = 16'b1010101000001000;
				18'b001110010100011100: oled_data = 16'b1011101001001001;
				18'b001110010110011100: oled_data = 16'b1011001001001001;
				18'b001110011000011100: oled_data = 16'b1010000111101000;
				18'b001110011010011100: oled_data = 16'b1010000111000111;
				18'b001110011100011100: oled_data = 16'b1011001001001001;
				18'b001110011110011100: oled_data = 16'b1011001000101000;
				18'b001110100000011100: oled_data = 16'b1011001000101001;
				18'b001110100010011100: oled_data = 16'b1011001000101000;
				18'b001110100100011100: oled_data = 16'b1011001000101000;
				18'b001110100110011100: oled_data = 16'b1010101000101000;
				18'b001100011000011101: oled_data = 16'b1101110011010110;
				18'b001100011010011101: oled_data = 16'b1010110000101010;
				18'b001100011100011101: oled_data = 16'b1011110001101110;
				18'b001100011110011101: oled_data = 16'b1101110011010110;
				18'b001100100000011101: oled_data = 16'b1101110011010110;
				18'b001100100010011101: oled_data = 16'b1100010000010011;
				18'b001100100100011101: oled_data = 16'b1100001111110010;
				18'b001100100110011101: oled_data = 16'b1110010011010110;
				18'b001100101000011101: oled_data = 16'b1101110010110101;
				18'b001100101010011101: oled_data = 16'b1101010101110110;
				18'b001100101100011101: oled_data = 16'b1110111011111010;
				18'b001100101110011101: oled_data = 16'b1101011000111000;
				18'b001100110000011101: oled_data = 16'b1101010100010101;
				18'b001100110010011101: oled_data = 16'b1101110010110101;
				18'b001100110100011101: oled_data = 16'b1101010010010100;
				18'b001100110110011101: oled_data = 16'b1101110011010110;
				18'b001100111000011101: oled_data = 16'b1101110011010101;
				18'b001100111010011101: oled_data = 16'b1101110011010101;
				18'b001100111100011101: oled_data = 16'b1101110011010101;
				18'b001100111110011101: oled_data = 16'b1101110011010101;
				18'b001101000000011101: oled_data = 16'b1101110011010101;
				18'b001101000010011101: oled_data = 16'b1101110011010110;
				18'b001101000100011101: oled_data = 16'b1101010011010100;
				18'b001101000110011101: oled_data = 16'b1101010101110110;
				18'b001101001000011101: oled_data = 16'b1100110010110100;
				18'b001101001010011101: oled_data = 16'b1110010011010110;
				18'b001101001100011101: oled_data = 16'b1101110010110101;
				18'b001101001110011101: oled_data = 16'b1101010100010101;
				18'b001101010000011101: oled_data = 16'b1101010010110100;
				18'b001101010010011101: oled_data = 16'b1101110010110101;
				18'b001101010100011101: oled_data = 16'b1101110010110101;
				18'b001101010110011101: oled_data = 16'b1101110010110101;
				18'b001101011000011101: oled_data = 16'b1101010100110110;
				18'b001101011010011101: oled_data = 16'b1110111011011011;
				18'b001101011100011101: oled_data = 16'b1101110101110111;
				18'b001101011110011101: oled_data = 16'b1101110010110101;
				18'b001101100000011101: oled_data = 16'b1101110011010110;
				18'b001101100010011101: oled_data = 16'b1101010010010100;
				18'b001101100100011101: oled_data = 16'b1011001101110000;
				18'b001101100110011101: oled_data = 16'b1011001101110000;
				18'b001101101000011101: oled_data = 16'b1011101110110001;
				18'b001101101010011101: oled_data = 16'b1100110001010011;
				18'b001101101100011101: oled_data = 16'b1101110010110101;
				18'b001101101110011101: oled_data = 16'b1101110011010101;
				18'b001101110000011101: oled_data = 16'b1101010110010111;
				18'b001101110010011101: oled_data = 16'b1101111001111001;
				18'b001101110100011101: oled_data = 16'b1110011011011010;
				18'b001101110110011101: oled_data = 16'b1011110001010010;
				18'b001101111000011101: oled_data = 16'b1100101111110010;
				18'b001101111010011101: oled_data = 16'b1101010001010100;
				18'b001101111100011101: oled_data = 16'b1100110000010011;
				18'b001101111110011101: oled_data = 16'b1011101110010000;
				18'b001110000000011101: oled_data = 16'b1110010011110011;
				18'b001110000010011101: oled_data = 16'b1110010011010011;
				18'b001110000100011101: oled_data = 16'b1011101010001010;
				18'b001110000110011101: oled_data = 16'b1011001000101001;
				18'b001110001000011101: oled_data = 16'b1100001011101011;
				18'b001110001010011101: oled_data = 16'b1100001100101100;
				18'b001110001100011101: oled_data = 16'b1011001000101001;
				18'b001110001110011101: oled_data = 16'b1011101001001001;
				18'b001110010000011101: oled_data = 16'b1011001000101000;
				18'b001110010010011101: oled_data = 16'b1011001001001001;
				18'b001110010100011101: oled_data = 16'b1011101001001001;
				18'b001110010110011101: oled_data = 16'b1010001000001000;
				18'b001110011000011101: oled_data = 16'b1001000101100110;
				18'b001110011010011101: oled_data = 16'b1010101000001000;
				18'b001110011100011101: oled_data = 16'b1011001000101001;
				18'b001110011110011101: oled_data = 16'b1011001000101000;
				18'b001110100000011101: oled_data = 16'b1011001000101001;
				18'b001110100010011101: oled_data = 16'b1011001000101000;
				18'b001110100100011101: oled_data = 16'b1011001000101000;
				18'b001110100110011101: oled_data = 16'b1010101000101000;
				18'b001100011000011110: oled_data = 16'b1101110010110101;
				18'b001100011010011110: oled_data = 16'b1011010001001001;
				18'b001100011100011110: oled_data = 16'b1011010001101100;
				18'b001100011110011110: oled_data = 16'b1101110011010110;
				18'b001100100000011110: oled_data = 16'b1101110011010110;
				18'b001100100010011110: oled_data = 16'b1100110001010100;
				18'b001100100100011110: oled_data = 16'b1011101110110001;
				18'b001100100110011110: oled_data = 16'b1110010011010110;
				18'b001100101000011110: oled_data = 16'b1101110010110101;
				18'b001100101010011110: oled_data = 16'b1101010101110110;
				18'b001100101100011110: oled_data = 16'b1110111100011011;
				18'b001100101110011110: oled_data = 16'b1110011010111001;
				18'b001100110000011110: oled_data = 16'b1100110101010101;
				18'b001100110010011110: oled_data = 16'b1101110010110101;
				18'b001100110100011110: oled_data = 16'b1101010010010100;
				18'b001100110110011110: oled_data = 16'b1101110011010101;
				18'b001100111000011110: oled_data = 16'b1101110011010101;
				18'b001100111010011110: oled_data = 16'b1101110011010101;
				18'b001100111100011110: oled_data = 16'b1101110011010101;
				18'b001100111110011110: oled_data = 16'b1101110011010101;
				18'b001101000000011110: oled_data = 16'b1101110011010101;
				18'b001101000010011110: oled_data = 16'b1101110011010110;
				18'b001101000100011110: oled_data = 16'b1101110010110101;
				18'b001101000110011110: oled_data = 16'b1101110111010111;
				18'b001101001000011110: oled_data = 16'b1101010101110110;
				18'b001101001010011110: oled_data = 16'b1101110010110101;
				18'b001101001100011110: oled_data = 16'b1101110011010101;
				18'b001101001110011110: oled_data = 16'b1101010110010111;
				18'b001101010000011110: oled_data = 16'b1100010010110100;
				18'b001101010010011110: oled_data = 16'b1101010001110100;
				18'b001101010100011110: oled_data = 16'b1101110011010101;
				18'b001101010110011110: oled_data = 16'b1101110011010101;
				18'b001101011000011110: oled_data = 16'b1101010011010101;
				18'b001101011010011110: oled_data = 16'b1110011010011010;
				18'b001101011100011110: oled_data = 16'b1110111011011010;
				18'b001101011110011110: oled_data = 16'b1101010101010110;
				18'b001101100000011110: oled_data = 16'b1101110011010101;
				18'b001101100010011110: oled_data = 16'b1101110011110110;
				18'b001101100100011110: oled_data = 16'b1101010001010100;
				18'b001101100110011110: oled_data = 16'b1100110000110011;
				18'b001101101000011110: oled_data = 16'b1101110010110101;
				18'b001101101010011110: oled_data = 16'b1101110011010110;
				18'b001101101100011110: oled_data = 16'b1101110011010101;
				18'b001101101110011110: oled_data = 16'b1101110011010110;
				18'b001101110000011110: oled_data = 16'b1100110010110100;
				18'b001101110010011110: oled_data = 16'b1101110110110111;
				18'b001101110100011110: oled_data = 16'b1110111100111011;
				18'b001101110110011110: oled_data = 16'b1100110100110101;
				18'b001101111000011110: oled_data = 16'b1011101101010000;
				18'b001101111010011110: oled_data = 16'b1011101101110001;
				18'b001101111100011110: oled_data = 16'b1011001101110000;
				18'b001101111110011110: oled_data = 16'b1011101111110000;
				18'b001110000000011110: oled_data = 16'b1110110100110100;
				18'b001110000010011110: oled_data = 16'b1101001111110000;
				18'b001110000100011110: oled_data = 16'b1011001000101001;
				18'b001110000110011110: oled_data = 16'b1011101001001001;
				18'b001110001000011110: oled_data = 16'b1100001100001100;
				18'b001110001010011110: oled_data = 16'b1011101010001010;
				18'b001110001100011110: oled_data = 16'b1011001001001001;
				18'b001110001110011110: oled_data = 16'b1011001001001001;
				18'b001110010000011110: oled_data = 16'b1010101000101000;
				18'b001110010010011110: oled_data = 16'b1011001001001001;
				18'b001110010100011110: oled_data = 16'b1010101000101000;
				18'b001110010110011110: oled_data = 16'b1000100101100110;
				18'b001110011000011110: oled_data = 16'b1001100110100111;
				18'b001110011010011110: oled_data = 16'b1011101010001010;
				18'b001110011100011110: oled_data = 16'b1011101010101010;
				18'b001110011110011110: oled_data = 16'b1011001000101000;
				18'b001110100000011110: oled_data = 16'b1011001000101001;
				18'b001110100010011110: oled_data = 16'b1011001000101000;
				18'b001110100100011110: oled_data = 16'b1011001000101000;
				18'b001110100110011110: oled_data = 16'b1010101000101000;
				18'b001100011000011111: oled_data = 16'b1101010010010100;
				18'b001100011010011111: oled_data = 16'b1011010001101010;
				18'b001100011100011111: oled_data = 16'b1011010000101011;
				18'b001100011110011111: oled_data = 16'b1101110010110101;
				18'b001100100000011111: oled_data = 16'b1101110011010110;
				18'b001100100010011111: oled_data = 16'b1101010010010101;
				18'b001100100100011111: oled_data = 16'b1011001101110001;
				18'b001100100110011111: oled_data = 16'b1101110010010101;
				18'b001100101000011111: oled_data = 16'b1101110010110101;
				18'b001100101010011111: oled_data = 16'b1101010101110110;
				18'b001100101100011111: oled_data = 16'b1110111100011011;
				18'b001100101110011111: oled_data = 16'b1110111100011010;
				18'b001100110000011111: oled_data = 16'b1101111000011000;
				18'b001100110010011111: oled_data = 16'b1100110010010100;
				18'b001100110100011111: oled_data = 16'b1101110010110101;
				18'b001100110110011111: oled_data = 16'b1101010010010101;
				18'b001100111000011111: oled_data = 16'b1101110011010110;
				18'b001100111010011111: oled_data = 16'b1101110011010101;
				18'b001100111100011111: oled_data = 16'b1101110011010101;
				18'b001100111110011111: oled_data = 16'b1101110011010101;
				18'b001101000000011111: oled_data = 16'b1101110011010101;
				18'b001101000010011111: oled_data = 16'b1101110011010110;
				18'b001101000100011111: oled_data = 16'b1101110011010101;
				18'b001101000110011111: oled_data = 16'b1101010101110110;
				18'b001101001000011111: oled_data = 16'b1110011001111001;
				18'b001101001010011111: oled_data = 16'b1101010010010100;
				18'b001101001100011111: oled_data = 16'b1101010001110100;
				18'b001101001110011111: oled_data = 16'b1100110101010110;
				18'b001101010000011111: oled_data = 16'b1110011001011001;
				18'b001101010010011111: oled_data = 16'b1101010011010101;
				18'b001101010100011111: oled_data = 16'b1101110011010101;
				18'b001101010110011111: oled_data = 16'b1101110011010101;
				18'b001101011000011111: oled_data = 16'b1101110010110101;
				18'b001101011010011111: oled_data = 16'b1101110111111000;
				18'b001101011100011111: oled_data = 16'b1110111100011011;
				18'b001101011110011111: oled_data = 16'b1110111010111010;
				18'b001101100000011111: oled_data = 16'b1100010010110100;
				18'b001101100010011111: oled_data = 16'b1101110010110101;
				18'b001101100100011111: oled_data = 16'b1101110011010101;
				18'b001101100110011111: oled_data = 16'b1101010010010100;
				18'b001101101000011111: oled_data = 16'b1101010010010100;
				18'b001101101010011111: oled_data = 16'b1101110011010110;
				18'b001101101100011111: oled_data = 16'b1101110011010101;
				18'b001101101110011111: oled_data = 16'b1101110011010110;
				18'b001101110000011111: oled_data = 16'b1101110011010110;
				18'b001101110010011111: oled_data = 16'b1101010100010101;
				18'b001101110100011111: oled_data = 16'b1110111011011011;
				18'b001101110110011111: oled_data = 16'b1101110111011000;
				18'b001101111000011111: oled_data = 16'b1011101101110001;
				18'b001101111010011111: oled_data = 16'b1011101110010001;
				18'b001101111100011111: oled_data = 16'b1010101101001111;
				18'b001101111110011111: oled_data = 16'b1101010010010010;
				18'b001110000000011111: oled_data = 16'b1110110100010100;
				18'b001110000010011111: oled_data = 16'b1100001100001101;
				18'b001110000100011111: oled_data = 16'b1011001000101001;
				18'b001110000110011111: oled_data = 16'b1011101001001001;
				18'b001110001000011111: oled_data = 16'b1011101010001010;
				18'b001110001010011111: oled_data = 16'b1011001001001001;
				18'b001110001100011111: oled_data = 16'b1011001001001001;
				18'b001110001110011111: oled_data = 16'b1010101000101000;
				18'b001110010000011111: oled_data = 16'b1011001001001001;
				18'b001110010010011111: oled_data = 16'b1011001000101001;
				18'b001110010100011111: oled_data = 16'b1001000110000111;
				18'b001110010110011111: oled_data = 16'b1001000101100110;
				18'b001110011000011111: oled_data = 16'b1011001001001010;
				18'b001110011010011111: oled_data = 16'b1101001111101111;
				18'b001110011100011111: oled_data = 16'b1011101010001010;
				18'b001110011110011111: oled_data = 16'b1011001000101000;
				18'b001110100000011111: oled_data = 16'b1011001000101001;
				18'b001110100010011111: oled_data = 16'b1011001000101000;
				18'b001110100100011111: oled_data = 16'b1011001000101000;
				18'b001110100110011111: oled_data = 16'b1010101000101000;
				18'b001100011000100000: oled_data = 16'b1101010001110100;
				18'b001100011010100000: oled_data = 16'b1011010001101001;
				18'b001100011100100000: oled_data = 16'b1011010001001011;
				18'b001100011110100000: oled_data = 16'b1101010010010101;
				18'b001100100000100000: oled_data = 16'b1110010011010110;
				18'b001100100010100000: oled_data = 16'b1101110010110101;
				18'b001100100100100000: oled_data = 16'b1011001110010001;
				18'b001100100110100000: oled_data = 16'b1100110001010100;
				18'b001100101000100000: oled_data = 16'b1101110011010110;
				18'b001100101010100000: oled_data = 16'b1010110000110001;
				18'b001100101100100000: oled_data = 16'b1101111001111000;
				18'b001100101110100000: oled_data = 16'b1110111100111011;
				18'b001100110000100000: oled_data = 16'b1110111100011011;
				18'b001100110010100000: oled_data = 16'b1100110101010101;
				18'b001100110100100000: oled_data = 16'b1101010010010100;
				18'b001100110110100000: oled_data = 16'b1101010001110100;
				18'b001100111000100000: oled_data = 16'b1101110011010101;
				18'b001100111010100000: oled_data = 16'b1101110011010101;
				18'b001100111100100000: oled_data = 16'b1101110011010101;
				18'b001100111110100000: oled_data = 16'b1101110011010101;
				18'b001101000000100000: oled_data = 16'b1101110010110101;
				18'b001101000010100000: oled_data = 16'b1101110010110101;
				18'b001101000100100000: oled_data = 16'b1101110010110101;
				18'b001101000110100000: oled_data = 16'b1100110011010101;
				18'b001101001000100000: oled_data = 16'b1101111001111000;
				18'b001101001010100000: oled_data = 16'b1100110011110101;
				18'b001101001100100000: oled_data = 16'b1101110010110101;
				18'b001101001110100000: oled_data = 16'b1101010100110110;
				18'b001101010000100000: oled_data = 16'b1110111100011011;
				18'b001101010010100000: oled_data = 16'b1110011001111001;
				18'b001101010100100000: oled_data = 16'b1101010100010101;
				18'b001101010110100000: oled_data = 16'b1110010011110110;
				18'b001101011000100000: oled_data = 16'b1101010010110101;
				18'b001101011010100000: oled_data = 16'b1011110010110011;
				18'b001101011100100000: oled_data = 16'b1110111011111010;
				18'b001101011110100000: oled_data = 16'b1110111100111011;
				18'b001101100000100000: oled_data = 16'b1100110101110101;
				18'b001101100010100000: oled_data = 16'b1011001111010001;
				18'b001101100100100000: oled_data = 16'b1101010010010100;
				18'b001101100110100000: oled_data = 16'b1110010011010110;
				18'b001101101000100000: oled_data = 16'b1101010010010100;
				18'b001101101010100000: oled_data = 16'b1101010010010100;
				18'b001101101100100000: oled_data = 16'b1101110011010101;
				18'b001101101110100000: oled_data = 16'b1101110011010110;
				18'b001101110000100000: oled_data = 16'b1101110011010101;
				18'b001101110010100000: oled_data = 16'b1101010011010101;
				18'b001101110100100000: oled_data = 16'b1101010101110110;
				18'b001101110110100000: oled_data = 16'b1101110111011000;
				18'b001101111000100000: oled_data = 16'b1011101101110001;
				18'b001101111010100000: oled_data = 16'b1011101101010001;
				18'b001101111100100000: oled_data = 16'b1011001101110000;
				18'b001101111110100000: oled_data = 16'b1110010011010011;
				18'b001110000000100000: oled_data = 16'b1110010011010011;
				18'b001110000010100000: oled_data = 16'b1011001001101010;
				18'b001110000100100000: oled_data = 16'b1011001000101001;
				18'b001110000110100000: oled_data = 16'b1011001001001001;
				18'b001110001000100000: oled_data = 16'b1011001001001001;
				18'b001110001010100000: oled_data = 16'b1011001001001001;
				18'b001110001100100000: oled_data = 16'b1011001001001001;
				18'b001110001110100000: oled_data = 16'b1010101000101001;
				18'b001110010000100000: oled_data = 16'b1011001001001001;
				18'b001110010010100000: oled_data = 16'b1001100110100111;
				18'b001110010100100000: oled_data = 16'b1000100101000110;
				18'b001110010110100000: oled_data = 16'b1010000111001000;
				18'b001110011000100000: oled_data = 16'b1100101101001101;
				18'b001110011010100000: oled_data = 16'b1100001100001100;
				18'b001110011100100000: oled_data = 16'b1011001000101000;
				18'b001110011110100000: oled_data = 16'b1011001000101001;
				18'b001110100000100000: oled_data = 16'b1011001000101001;
				18'b001110100010100000: oled_data = 16'b1011001000101000;
				18'b001110100100100000: oled_data = 16'b1011001000101000;
				18'b001110100110100000: oled_data = 16'b1010101000101000;
				18'b001100011000100001: oled_data = 16'b1101010010110011;
				18'b001100011010100001: oled_data = 16'b1011110010001011;
				18'b001100011100100001: oled_data = 16'b1100010010010000;
				18'b001100011110100001: oled_data = 16'b1101010001010100;
				18'b001100100000100001: oled_data = 16'b1101110011010101;
				18'b001100100010100001: oled_data = 16'b1101110011010101;
				18'b001100100100100001: oled_data = 16'b1011101110110001;
				18'b001100100110100001: oled_data = 16'b1100001111110011;
				18'b001100101000100001: oled_data = 16'b1110010100010110;
				18'b001100101010100001: oled_data = 16'b1000001011001100;
				18'b001100101100100001: oled_data = 16'b0101101001001000;
				18'b001100101110100001: oled_data = 16'b1100111000110111;
				18'b001100110000100001: oled_data = 16'b1110111100111011;
				18'b001100110010100001: oled_data = 16'b1110011010111001;
				18'b001100110100100001: oled_data = 16'b1100110010110100;
				18'b001100110110100001: oled_data = 16'b1101110010010100;
				18'b001100111000100001: oled_data = 16'b1101110010010101;
				18'b001100111010100001: oled_data = 16'b1101110011010110;
				18'b001100111100100001: oled_data = 16'b1101110011010101;
				18'b001100111110100001: oled_data = 16'b1101010010010100;
				18'b001101000000100001: oled_data = 16'b1100110001010011;
				18'b001101000010100001: oled_data = 16'b1101010001010100;
				18'b001101000100100001: oled_data = 16'b1101010001110100;
				18'b001101000110100001: oled_data = 16'b1101010011010100;
				18'b001101001000100001: oled_data = 16'b1110011010111010;
				18'b001101001010100001: oled_data = 16'b1110011000111001;
				18'b001101001100100001: oled_data = 16'b1101110011010101;
				18'b001101001110100001: oled_data = 16'b1101010100010101;
				18'b001101010000100001: oled_data = 16'b1110011011011010;
				18'b001101010010100001: oled_data = 16'b1110111101011100;
				18'b001101010100100001: oled_data = 16'b1101111000111001;
				18'b001101010110100001: oled_data = 16'b1001101111010000;
				18'b001101011000100001: oled_data = 16'b0111001000101010;
				18'b001101011010100001: oled_data = 16'b1000101100001101;
				18'b001101011100100001: oled_data = 16'b1110011010011001;
				18'b001101011110100001: oled_data = 16'b1110111100111010;
				18'b001101100000100001: oled_data = 16'b1110011010111001;
				18'b001101100010100001: oled_data = 16'b1010101110110000;
				18'b001101100100100001: oled_data = 16'b1011001101110000;
				18'b001101100110100001: oled_data = 16'b1100001111110010;
				18'b001101101000100001: oled_data = 16'b1101010010010101;
				18'b001101101010100001: oled_data = 16'b1101010010010101;
				18'b001101101100100001: oled_data = 16'b1101010001110100;
				18'b001101101110100001: oled_data = 16'b1101010001110100;
				18'b001101110000100001: oled_data = 16'b1101010010010100;
				18'b001101110010100001: oled_data = 16'b1101110011010101;
				18'b001101110100100001: oled_data = 16'b1101010011010101;
				18'b001101110110100001: oled_data = 16'b1100110011010101;
				18'b001101111000100001: oled_data = 16'b1011101110010001;
				18'b001101111010100001: oled_data = 16'b1010101100001111;
				18'b001101111100100001: oled_data = 16'b1011101110110000;
				18'b001101111110100001: oled_data = 16'b1110010100010100;
				18'b001110000000100001: oled_data = 16'b1101110001110001;
				18'b001110000010100001: oled_data = 16'b1011001000101001;
				18'b001110000100100001: oled_data = 16'b1011001001001001;
				18'b001110000110100001: oled_data = 16'b1011001001001001;
				18'b001110001000100001: oled_data = 16'b1011001001001001;
				18'b001110001010100001: oled_data = 16'b1011001001001001;
				18'b001110001100100001: oled_data = 16'b1010101000101001;
				18'b001110001110100001: oled_data = 16'b1011001001001001;
				18'b001110010000100001: oled_data = 16'b1010000111101000;
				18'b001110010010100001: oled_data = 16'b1000100101000110;
				18'b001110010100100001: oled_data = 16'b1001100110000111;
				18'b001110010110100001: oled_data = 16'b1011001000101001;
				18'b001110011000100001: oled_data = 16'b1011101010001010;
				18'b001110011010100001: oled_data = 16'b1011001001001001;
				18'b001110011100100001: oled_data = 16'b1011001000101001;
				18'b001110011110100001: oled_data = 16'b1011001000101001;
				18'b001110100000100001: oled_data = 16'b1011001000101001;
				18'b001110100010100001: oled_data = 16'b1011001000101000;
				18'b001110100100100001: oled_data = 16'b1011001000101000;
				18'b001110100110100001: oled_data = 16'b1010101000101000;
				18'b001100011000100010: oled_data = 16'b1011010000110000;
				18'b001100011010100010: oled_data = 16'b1011010000001101;
				18'b001100011100100010: oled_data = 16'b1101110010110101;
				18'b001100011110100010: oled_data = 16'b1101010001010011;
				18'b001100100000100010: oled_data = 16'b1101010010010101;
				18'b001100100010100010: oled_data = 16'b1101110011110110;
				18'b001100100100100010: oled_data = 16'b1100001111010010;
				18'b001100100110100010: oled_data = 16'b1011001101110001;
				18'b001100101000100010: oled_data = 16'b1101110011010110;
				18'b001100101010100010: oled_data = 16'b1011001111010001;
				18'b001100101100100010: oled_data = 16'b0011000100000100;
				18'b001100101110100010: oled_data = 16'b0100101000000111;
				18'b001100110000100010: oled_data = 16'b1100111000110111;
				18'b001100110010100010: oled_data = 16'b1111011101011011;
				18'b001100110100100010: oled_data = 16'b1101010111010111;
				18'b001100110110100010: oled_data = 16'b1101110010110101;
				18'b001100111000100010: oled_data = 16'b1101010001110100;
				18'b001100111010100010: oled_data = 16'b1101110011010101;
				18'b001100111100100010: oled_data = 16'b1101110011010101;
				18'b001100111110100010: oled_data = 16'b1101110011010110;
				18'b001101000000100010: oled_data = 16'b1101110011010110;
				18'b001101000010100010: oled_data = 16'b1110010011010110;
				18'b001101000100100010: oled_data = 16'b1110010011010110;
				18'b001101000110100010: oled_data = 16'b1101110011010101;
				18'b001101001000100010: oled_data = 16'b1110011010011001;
				18'b001101001010100010: oled_data = 16'b1110011011011010;
				18'b001101001100100010: oled_data = 16'b1101010100010101;
				18'b001101001110100010: oled_data = 16'b1101110011110101;
				18'b001101010000100010: oled_data = 16'b1110011001111001;
				18'b001101010010100010: oled_data = 16'b1011110110110101;
				18'b001101010100100010: oled_data = 16'b0110001011001011;
				18'b001101010110100010: oled_data = 16'b0011000101000100;
				18'b001101011000100010: oled_data = 16'b0101101000001000;
				18'b001101011010100010: oled_data = 16'b1010101111010000;
				18'b001101011100100010: oled_data = 16'b1101110111010111;
				18'b001101011110100010: oled_data = 16'b1110111100011010;
				18'b001101100000100010: oled_data = 16'b1110111100111011;
				18'b001101100010100010: oled_data = 16'b1100010100010100;
				18'b001101100100100010: oled_data = 16'b1011001101010000;
				18'b001101100110100010: oled_data = 16'b1011001101110001;
				18'b001101101000100010: oled_data = 16'b1011001101110001;
				18'b001101101010100010: oled_data = 16'b1011101110110010;
				18'b001101101100100010: oled_data = 16'b1100001111110011;
				18'b001101101110100010: oled_data = 16'b1100010000010011;
				18'b001101110000100010: oled_data = 16'b1100110001010011;
				18'b001101110010100010: oled_data = 16'b1101110011110101;
				18'b001101110100100010: oled_data = 16'b1101110011010101;
				18'b001101110110100010: oled_data = 16'b1101110010110101;
				18'b001101111000100010: oled_data = 16'b1100010000010010;
				18'b001101111010100010: oled_data = 16'b1011001110010001;
				18'b001101111100100010: oled_data = 16'b1100001111110001;
				18'b001101111110100010: oled_data = 16'b1110110100110101;
				18'b001110000000100010: oled_data = 16'b1100101111001111;
				18'b001110000010100010: oled_data = 16'b1010101000001000;
				18'b001110000100100010: oled_data = 16'b1011101001001001;
				18'b001110000110100010: oled_data = 16'b1011001001001001;
				18'b001110001000100010: oled_data = 16'b1011001001001001;
				18'b001110001010100010: oled_data = 16'b1011001001001001;
				18'b001110001100100010: oled_data = 16'b1010101000101000;
				18'b001110001110100010: oled_data = 16'b1011001001001001;
				18'b001110010000100010: oled_data = 16'b1001000101100111;
				18'b001110010010100010: oled_data = 16'b1000100101000110;
				18'b001110010100100010: oled_data = 16'b1010101000001000;
				18'b001110010110100010: oled_data = 16'b1011001001001001;
				18'b001110011000100010: oled_data = 16'b1011001001001001;
				18'b001110011010100010: oled_data = 16'b1011001001001001;
				18'b001110011100100010: oled_data = 16'b1011001001001001;
				18'b001110011110100010: oled_data = 16'b1011001001001001;
				18'b001110100000100010: oled_data = 16'b1011001000101001;
				18'b001110100010100010: oled_data = 16'b1011001000101000;
				18'b001110100100100010: oled_data = 16'b1011001000001000;
				18'b001110100110100010: oled_data = 16'b1010101000001000;
				18'b001100011000100011: oled_data = 16'b0111001001101011;
				18'b001100011010100011: oled_data = 16'b1010001110001111;
				18'b001100011100100011: oled_data = 16'b1101110011010101;
				18'b001100011110100011: oled_data = 16'b1101010010010100;
				18'b001100100000100011: oled_data = 16'b1100001111110010;
				18'b001100100010100011: oled_data = 16'b1110010011110110;
				18'b001100100100100011: oled_data = 16'b1100110000110011;
				18'b001100100110100011: oled_data = 16'b1011001101110001;
				18'b001100101000100011: oled_data = 16'b1100110001010100;
				18'b001100101010100011: oled_data = 16'b1101110100110110;
				18'b001100101100100011: oled_data = 16'b1010010010110010;
				18'b001100101110100011: oled_data = 16'b0011100101100100;
				18'b001100110000100011: oled_data = 16'b0101001001001000;
				18'b001100110010100011: oled_data = 16'b1101011001111000;
				18'b001100110100100011: oled_data = 16'b1110111100011010;
				18'b001100110110100011: oled_data = 16'b1101010100110101;
				18'b001100111000100011: oled_data = 16'b1101010010010100;
				18'b001100111010100011: oled_data = 16'b1101110010010101;
				18'b001100111100100011: oled_data = 16'b1110010011010110;
				18'b001100111110100011: oled_data = 16'b1101110011010101;
				18'b001101000000100011: oled_data = 16'b1101110011010101;
				18'b001101000010100011: oled_data = 16'b1101110011010101;
				18'b001101000100100011: oled_data = 16'b1110010010110101;
				18'b001101000110100011: oled_data = 16'b1101010011010101;
				18'b001101001000100011: oled_data = 16'b1110011001111001;
				18'b001101001010100011: oled_data = 16'b1110111100111011;
				18'b001101001100100011: oled_data = 16'b1101111000011000;
				18'b001101001110100011: oled_data = 16'b1100010001110011;
				18'b001101010000100011: oled_data = 16'b0111101100001100;
				18'b001101010010100011: oled_data = 16'b0011000101000100;
				18'b001101010100100011: oled_data = 16'b0011100110000110;
				18'b001101010110100011: oled_data = 16'b1000110000110000;
				18'b001101011000100011: oled_data = 16'b1101011000011000;
				18'b001101011010100011: oled_data = 16'b1101010100010101;
				18'b001101011100100011: oled_data = 16'b1101010011110101;
				18'b001101011110100011: oled_data = 16'b1110011010111010;
				18'b001101100000100011: oled_data = 16'b1110111100111011;
				18'b001101100010100011: oled_data = 16'b1110011010011001;
				18'b001101100100100011: oled_data = 16'b1011001111110001;
				18'b001101100110100011: oled_data = 16'b1011101111010010;
				18'b001101101000100011: oled_data = 16'b1100110001110100;
				18'b001101101010100011: oled_data = 16'b1100110001110100;
				18'b001101101100100011: oled_data = 16'b1101010001110101;
				18'b001101101110100011: oled_data = 16'b1101010010110101;
				18'b001101110000100011: oled_data = 16'b1101010010110101;
				18'b001101110010100011: oled_data = 16'b1101110011010101;
				18'b001101110100100011: oled_data = 16'b1101110011010101;
				18'b001101110110100011: oled_data = 16'b1101110011010101;
				18'b001101111000100011: oled_data = 16'b1100110001010011;
				18'b001101111010100011: oled_data = 16'b1100110001010011;
				18'b001101111100100011: oled_data = 16'b1101010001110011;
				18'b001101111110100011: oled_data = 16'b1110110100010100;
				18'b001110000000100011: oled_data = 16'b1100001100101100;
				18'b001110000010100011: oled_data = 16'b1010101000101000;
				18'b001110000100100011: oled_data = 16'b1011101001001001;
				18'b001110000110100011: oled_data = 16'b1011001001001001;
				18'b001110001000100011: oled_data = 16'b1011001001001001;
				18'b001110001010100011: oled_data = 16'b1011001000101001;
				18'b001110001100100011: oled_data = 16'b1010101000101001;
				18'b001110001110100011: oled_data = 16'b1010000111101000;
				18'b001110010000100011: oled_data = 16'b1000100101000110;
				18'b001110010010100011: oled_data = 16'b1001100111001000;
				18'b001110010100100011: oled_data = 16'b1011001001001001;
				18'b001110010110100011: oled_data = 16'b1011001001001001;
				18'b001110011000100011: oled_data = 16'b1011001001001001;
				18'b001110011010100011: oled_data = 16'b1011001001001001;
				18'b001110011100100011: oled_data = 16'b1011001000101001;
				18'b001110011110100011: oled_data = 16'b1011001000101001;
				18'b001110100000100011: oled_data = 16'b1011001000101001;
				18'b001110100010100011: oled_data = 16'b1011001000101000;
				18'b001110100100100011: oled_data = 16'b1011001000001000;
				18'b001110100110100011: oled_data = 16'b1010101000001000;
				18'b001100011000100100: oled_data = 16'b0100000111000111;
				18'b001100011010100100: oled_data = 16'b1010101111110001;
				18'b001100011100100100: oled_data = 16'b1110010011110110;
				18'b001100011110100100: oled_data = 16'b1101110011010101;
				18'b001100100000100100: oled_data = 16'b1011101110010001;
				18'b001100100010100100: oled_data = 16'b1100110001010011;
				18'b001100100100100100: oled_data = 16'b1101010001110100;
				18'b001100100110100100: oled_data = 16'b1011001101110001;
				18'b001100101000100100: oled_data = 16'b1011001110110010;
				18'b001100101010100100: oled_data = 16'b1101010010110101;
				18'b001100101100100100: oled_data = 16'b1110111010011010;
				18'b001100101110100100: oled_data = 16'b1011110110110101;
				18'b001100110000100100: oled_data = 16'b0100101000000111;
				18'b001100110010100100: oled_data = 16'b0110001011001010;
				18'b001100110100100100: oled_data = 16'b1110011011011010;
				18'b001100110110100100: oled_data = 16'b1110011010111001;
				18'b001100111000100100: oled_data = 16'b1101010011110101;
				18'b001100111010100100: oled_data = 16'b1101010001010100;
				18'b001100111100100100: oled_data = 16'b1101110010110101;
				18'b001100111110100100: oled_data = 16'b1110010011010101;
				18'b001101000000100100: oled_data = 16'b1101110011010101;
				18'b001101000010100100: oled_data = 16'b1101110011010101;
				18'b001101000100100100: oled_data = 16'b1110010011010101;
				18'b001101000110100100: oled_data = 16'b1101110010110101;
				18'b001101001000100100: oled_data = 16'b1110011001111001;
				18'b001101001010100100: oled_data = 16'b1110111011111010;
				18'b001101001100100100: oled_data = 16'b1001110001110001;
				18'b001101001110100100: oled_data = 16'b0101000111101000;
				18'b001101010000100100: oled_data = 16'b0011100100100100;
				18'b001101010010100100: oled_data = 16'b0110001011001011;
				18'b001101010100100100: oled_data = 16'b1100110111110111;
				18'b001101010110100100: oled_data = 16'b1110111101011011;
				18'b001101011000100100: oled_data = 16'b1110111100111011;
				18'b001101011010100100: oled_data = 16'b1110011010111010;
				18'b001101011100100100: oled_data = 16'b1101010101110110;
				18'b001101011110100100: oled_data = 16'b1101010111010111;
				18'b001101100000100100: oled_data = 16'b1110111100011010;
				18'b001101100010100100: oled_data = 16'b1110111100111011;
				18'b001101100100100100: oled_data = 16'b1100110110010110;
				18'b001101100110100100: oled_data = 16'b1011001110110000;
				18'b001101101000100100: oled_data = 16'b1101110010010101;
				18'b001101101010100100: oled_data = 16'b1101110011010110;
				18'b001101101100100100: oled_data = 16'b1110010011010110;
				18'b001101101110100100: oled_data = 16'b1101110011010110;
				18'b001101110000100100: oled_data = 16'b1101110011010110;
				18'b001101110010100100: oled_data = 16'b1101110011010101;
				18'b001101110100100100: oled_data = 16'b1101110011010110;
				18'b001101110110100100: oled_data = 16'b1101010001110100;
				18'b001101111000100100: oled_data = 16'b1101110010110101;
				18'b001101111010100100: oled_data = 16'b1101110011010101;
				18'b001101111100100100: oled_data = 16'b1101010010110011;
				18'b001101111110100100: oled_data = 16'b1110110011110011;
				18'b001110000000100100: oled_data = 16'b1011001010101011;
				18'b001110000010100100: oled_data = 16'b1011001000101001;
				18'b001110000100100100: oled_data = 16'b1011001001001001;
				18'b001110000110100100: oled_data = 16'b1011001001001001;
				18'b001110001000100100: oled_data = 16'b1011001001001001;
				18'b001110001010100100: oled_data = 16'b1010101000101000;
				18'b001110001100100100: oled_data = 16'b1011001000101001;
				18'b001110001110100100: oled_data = 16'b1001000101100110;
				18'b001110010000100100: oled_data = 16'b1001000101100111;
				18'b001110010010100100: oled_data = 16'b1011001000101001;
				18'b001110010100100100: oled_data = 16'b1011001001001001;
				18'b001110010110100100: oled_data = 16'b1011001001101010;
				18'b001110011000100100: oled_data = 16'b1011001001001001;
				18'b001110011010100100: oled_data = 16'b1011001000101001;
				18'b001110011100100100: oled_data = 16'b1011001001001001;
				18'b001110011110100100: oled_data = 16'b1011001001001001;
				18'b001110100000100100: oled_data = 16'b1011001000101001;
				18'b001110100010100100: oled_data = 16'b1011001000101000;
				18'b001110100100100100: oled_data = 16'b1010101000101000;
				18'b001110100110100100: oled_data = 16'b1010101000101000;
				18'b001100011000100101: oled_data = 16'b0100000110100110;
				18'b001100011010100101: oled_data = 16'b1001101101001111;
				18'b001100011100100101: oled_data = 16'b1101110010110110;
				18'b001100011110100101: oled_data = 16'b1101110011010110;
				18'b001100100000100101: oled_data = 16'b1100110000010011;
				18'b001100100010100101: oled_data = 16'b1011001101110000;
				18'b001100100100100101: oled_data = 16'b1101010001110100;
				18'b001100100110100101: oled_data = 16'b1011101110010001;
				18'b001100101000100101: oled_data = 16'b1011110000110011;
				18'b001100101010100101: oled_data = 16'b1100110100010110;
				18'b001100101100100101: oled_data = 16'b1101111000011000;
				18'b001100101110100101: oled_data = 16'b1111011101111011;
				18'b001100110000100101: oled_data = 16'b1100111000010111;
				18'b001100110010100101: oled_data = 16'b0100100111100111;
				18'b001100110100100101: oled_data = 16'b0111001100101100;
				18'b001100110110100101: oled_data = 16'b1110111100011011;
				18'b001100111000100101: oled_data = 16'b1101111001111001;
				18'b001100111010100101: oled_data = 16'b1101010011010100;
				18'b001100111100100101: oled_data = 16'b1101010001110100;
				18'b001100111110100101: oled_data = 16'b1110010011010110;
				18'b001101000000100101: oled_data = 16'b1110010011010101;
				18'b001101000010100101: oled_data = 16'b1110010011010101;
				18'b001101000100100101: oled_data = 16'b1110010010110101;
				18'b001101000110100101: oled_data = 16'b1110010011110110;
				18'b001101001000100101: oled_data = 16'b1100110101110110;
				18'b001101001010100101: oled_data = 16'b0110101011001011;
				18'b001101001100100101: oled_data = 16'b0011000100100100;
				18'b001101001110100101: oled_data = 16'b0100100111100111;
				18'b001101010000100101: oled_data = 16'b1001110001010000;
				18'b001101010010100101: oled_data = 16'b1110111100011011;
				18'b001101010100100101: oled_data = 16'b1110111100111011;
				18'b001101010110100101: oled_data = 16'b1110111100011010;
				18'b001101011000100101: oled_data = 16'b1110111100011010;
				18'b001101011010100101: oled_data = 16'b1110111100011011;
				18'b001101011100100101: oled_data = 16'b1110111100011011;
				18'b001101011110100101: oled_data = 16'b1110011010011001;
				18'b001101100000100101: oled_data = 16'b1110011100011010;
				18'b001101100010100101: oled_data = 16'b1110111100011011;
				18'b001101100100100101: oled_data = 16'b1110111011111010;
				18'b001101100110100101: oled_data = 16'b1011110001110010;
				18'b001101101000100101: oled_data = 16'b1100101111110010;
				18'b001101101010100101: oled_data = 16'b1110010010110110;
				18'b001101101100100101: oled_data = 16'b1110010010110110;
				18'b001101101110100101: oled_data = 16'b1110010010110110;
				18'b001101110000100101: oled_data = 16'b1110010010110110;
				18'b001101110010100101: oled_data = 16'b1101110011010110;
				18'b001101110100100101: oled_data = 16'b1101010010010101;
				18'b001101110110100101: oled_data = 16'b1101010001110100;
				18'b001101111000100101: oled_data = 16'b1101110011010101;
				18'b001101111010100101: oled_data = 16'b1101110010110101;
				18'b001101111100100101: oled_data = 16'b1101010010110011;
				18'b001101111110100101: oled_data = 16'b1110010011010011;
				18'b001110000000100101: oled_data = 16'b1010101001101001;
				18'b001110000010100101: oled_data = 16'b1011001001001001;
				18'b001110000100100101: oled_data = 16'b1011001001001001;
				18'b001110000110100101: oled_data = 16'b1011001001001001;
				18'b001110001000100101: oled_data = 16'b1011101010101010;
				18'b001110001010100101: oled_data = 16'b1011001010001001;
				18'b001110001100100101: oled_data = 16'b1010000111100111;
				18'b001110001110100101: oled_data = 16'b1000100101000110;
				18'b001110010000100101: oled_data = 16'b1010000111101001;
				18'b001110010010100101: oled_data = 16'b1011001001001001;
				18'b001110010100100101: oled_data = 16'b1011001000001001;
				18'b001110010110100101: oled_data = 16'b1011110010010010;
				18'b001110011000100101: oled_data = 16'b1011001011101100;
				18'b001110011010100101: oled_data = 16'b1011001000101001;
				18'b001110011100100101: oled_data = 16'b1011101010001010;
				18'b001110011110100101: oled_data = 16'b1011001001001001;
				18'b001110100000100101: oled_data = 16'b1011001000101001;
				18'b001110100010100101: oled_data = 16'b1011001000101000;
				18'b001110100100100101: oled_data = 16'b1010101000101000;
				18'b001110100110100101: oled_data = 16'b1010101000101000;
				18'b001100011000100110: oled_data = 16'b0100000111100111;
				18'b001100011010100110: oled_data = 16'b1011110000110010;
				18'b001100011100100110: oled_data = 16'b1100110000110011;
				18'b001100011110100110: oled_data = 16'b1101110011110110;
				18'b001100100000100110: oled_data = 16'b1101110010110101;
				18'b001100100010100110: oled_data = 16'b1011101110110001;
				18'b001100100100100110: oled_data = 16'b1011001110010000;
				18'b001100100110100110: oled_data = 16'b1011001101110001;
				18'b001100101000100110: oled_data = 16'b1011110001110100;
				18'b001100101010100110: oled_data = 16'b1101011000011000;
				18'b001100101100100110: oled_data = 16'b1100110110110110;
				18'b001100101110100110: oled_data = 16'b1110111100111011;
				18'b001100110000100110: oled_data = 16'b1111011101111100;
				18'b001100110010100110: oled_data = 16'b1100111000111000;
				18'b001100110100100110: oled_data = 16'b0100000111100111;
				18'b001100110110100110: oled_data = 16'b1001010001110000;
				18'b001100111000100110: oled_data = 16'b1111011101011011;
				18'b001100111010100110: oled_data = 16'b1101110111110111;
				18'b001100111100100110: oled_data = 16'b1100110001110100;
				18'b001100111110100110: oled_data = 16'b1101110010010101;
				18'b001101000000100110: oled_data = 16'b1101110011010110;
				18'b001101000010100110: oled_data = 16'b1101110011010101;
				18'b001101000100100110: oled_data = 16'b1110010011010110;
				18'b001101000110100110: oled_data = 16'b1100010000110011;
				18'b001101001000100110: oled_data = 16'b0101000111000111;
				18'b001101001010100110: oled_data = 16'b0011000101100101;
				18'b001101001100100110: oled_data = 16'b0111101110101110;
				18'b001101001110100110: oled_data = 16'b1100010101010101;
				18'b001101010000100110: oled_data = 16'b1101010110110110;
				18'b001101010010100110: oled_data = 16'b1110111100111011;
				18'b001101010100100110: oled_data = 16'b1110111100011010;
				18'b001101010110100110: oled_data = 16'b1110111100011010;
				18'b001101011000100110: oled_data = 16'b1110111100011010;
				18'b001101011010100110: oled_data = 16'b1110111100011010;
				18'b001101011100100110: oled_data = 16'b1110111100011011;
				18'b001101011110100110: oled_data = 16'b1110111100011011;
				18'b001101100000100110: oled_data = 16'b1110111100011010;
				18'b001101100010100110: oled_data = 16'b1110111100011010;
				18'b001101100100100110: oled_data = 16'b1110111100111011;
				18'b001101100110100110: oled_data = 16'b1110011001111001;
				18'b001101101000100110: oled_data = 16'b1011101111110001;
				18'b001101101010100110: oled_data = 16'b1101010001110100;
				18'b001101101100100110: oled_data = 16'b1110010011010101;
				18'b001101101110100110: oled_data = 16'b1101110010110101;
				18'b001101110000100110: oled_data = 16'b1101010001110101;
				18'b001101110010100110: oled_data = 16'b1101110010110101;
				18'b001101110100100110: oled_data = 16'b1101010001110100;
				18'b001101110110100110: oled_data = 16'b1101110010110101;
				18'b001101111000100110: oled_data = 16'b1101110011010101;
				18'b001101111010100110: oled_data = 16'b1101010010110101;
				18'b001101111100100110: oled_data = 16'b1101110011010100;
				18'b001101111110100110: oled_data = 16'b1101110001110001;
				18'b001110000000100110: oled_data = 16'b1010101000101001;
				18'b001110000010100110: oled_data = 16'b1011001001001001;
				18'b001110000100100110: oled_data = 16'b1011001010101010;
				18'b001110000110100110: oled_data = 16'b1101010000110000;
				18'b001110001000100110: oled_data = 16'b1110010010110011;
				18'b001110001010100110: oled_data = 16'b1100101110101111;
				18'b001110001100100110: oled_data = 16'b1010000111101000;
				18'b001110001110100110: oled_data = 16'b1001100110000111;
				18'b001110010000100110: oled_data = 16'b1011001001101010;
				18'b001110010010100110: oled_data = 16'b1011001001001001;
				18'b001110010100100110: oled_data = 16'b1011001010101011;
				18'b001110010110100110: oled_data = 16'b1100011010011010;
				18'b001110011000100110: oled_data = 16'b1011010010010010;
				18'b001110011010100110: oled_data = 16'b1011001000001000;
				18'b001110011100100110: oled_data = 16'b1011001000101001;
				18'b001110011110100110: oled_data = 16'b1011001000101001;
				18'b001110100000100110: oled_data = 16'b1011001000101001;
				18'b001110100010100110: oled_data = 16'b1011001000101000;
				18'b001110100100100110: oled_data = 16'b1010101000101000;
				18'b001110100110100110: oled_data = 16'b1010101000101000;
				18'b001100011000100111: oled_data = 16'b0011100111000110;
				18'b001100011010100111: oled_data = 16'b1100110010010100;
				18'b001100011100100111: oled_data = 16'b1101110010110101;
				18'b001100011110100111: oled_data = 16'b1101110011010110;
				18'b001100100000100111: oled_data = 16'b1110010011010110;
				18'b001100100010100111: oled_data = 16'b1100110000010011;
				18'b001100100100100111: oled_data = 16'b1010101100001111;
				18'b001100100110100111: oled_data = 16'b1010101100110000;
				18'b001100101000100111: oled_data = 16'b1011110001110100;
				18'b001100101010100111: oled_data = 16'b1110111100011011;
				18'b001100101100100111: oled_data = 16'b1100110111010110;
				18'b001100101110100111: oled_data = 16'b1101011010011000;
				18'b001100110000100111: oled_data = 16'b1100010111010110;
				18'b001100110010100111: oled_data = 16'b1010110100110100;
				18'b001100110100100111: oled_data = 16'b0110001010101011;
				18'b001100110110100111: oled_data = 16'b0011100110100110;
				18'b001100111000100111: oled_data = 16'b1101111010011001;
				18'b001100111010100111: oled_data = 16'b1110111100011011;
				18'b001100111100100111: oled_data = 16'b1101010111010111;
				18'b001100111110100111: oled_data = 16'b1100010001110011;
				18'b001101000000100111: oled_data = 16'b1101110010110101;
				18'b001101000010100111: oled_data = 16'b1101110011010110;
				18'b001101000100100111: oled_data = 16'b1110010011110110;
				18'b001101000110100111: oled_data = 16'b1000101010101100;
				18'b001101001000100111: oled_data = 16'b0011000100000100;
				18'b001101001010100111: oled_data = 16'b0101101010101010;
				18'b001101001100100111: oled_data = 16'b1100111000011000;
				18'b001101001110100111: oled_data = 16'b1101111001011001;
				18'b001101010000100111: oled_data = 16'b1101010110110110;
				18'b001101010010100111: oled_data = 16'b1111011101011100;
				18'b001101010100100111: oled_data = 16'b1110111100111011;
				18'b001101010110100111: oled_data = 16'b1110111100011011;
				18'b001101011000100111: oled_data = 16'b1110111100011011;
				18'b001101011010100111: oled_data = 16'b1110111100011011;
				18'b001101011100100111: oled_data = 16'b1110111100011011;
				18'b001101011110100111: oled_data = 16'b1110111100011011;
				18'b001101100000100111: oled_data = 16'b1110111100011011;
				18'b001101100010100111: oled_data = 16'b1110111100011010;
				18'b001101100100100111: oled_data = 16'b1110111100011010;
				18'b001101100110100111: oled_data = 16'b1110111100111011;
				18'b001101101000100111: oled_data = 16'b1101011000011000;
				18'b001101101010100111: oled_data = 16'b1011110000010010;
				18'b001101101100100111: oled_data = 16'b1101110010110101;
				18'b001101101110100111: oled_data = 16'b1101110011010101;
				18'b001101110000100111: oled_data = 16'b1101010010010101;
				18'b001101110010100111: oled_data = 16'b1100110000110011;
				18'b001101110100100111: oled_data = 16'b1101110011010101;
				18'b001101110110100111: oled_data = 16'b1101110011010101;
				18'b001101111000100111: oled_data = 16'b1101110011010101;
				18'b001101111010100111: oled_data = 16'b1101010010110101;
				18'b001101111100100111: oled_data = 16'b1101110011010100;
				18'b001101111110100111: oled_data = 16'b1101010000110000;
				18'b001110000000100111: oled_data = 16'b1010101000101000;
				18'b001110000010100111: oled_data = 16'b1011001001001001;
				18'b001110000100100111: oled_data = 16'b1101010001010001;
				18'b001110000110100111: oled_data = 16'b1110110011110011;
				18'b001110001000100111: oled_data = 16'b1100001100001101;
				18'b001110001010100111: oled_data = 16'b1011001000101001;
				18'b001110001100100111: oled_data = 16'b1011001000101001;
				18'b001110001110100111: oled_data = 16'b1011001001001001;
				18'b001110010000100111: oled_data = 16'b1011001001101010;
				18'b001110010010100111: oled_data = 16'b1011001000101001;
				18'b001110010100100111: oled_data = 16'b1011110001110010;
				18'b001110010110100111: oled_data = 16'b1011111100111100;
				18'b001110011000100111: oled_data = 16'b1011111000111000;
				18'b001110011010100111: oled_data = 16'b1011001001101010;
				18'b001110011100100111: oled_data = 16'b1011001000101001;
				18'b001110011110100111: oled_data = 16'b1011001001001001;
				18'b001110100000100111: oled_data = 16'b1011001000101000;
				18'b001110100010100111: oled_data = 16'b1010101000001000;
				18'b001110100100100111: oled_data = 16'b1010000111101000;
				18'b001110100110100111: oled_data = 16'b1010101000001000;
				18'b001100011000101000: oled_data = 16'b0101101001101001;
				18'b001100011010101000: oled_data = 16'b1101110010110101;
				18'b001100011100101000: oled_data = 16'b1110010011010110;
				18'b001100011110101000: oled_data = 16'b1101110011010110;
				18'b001100100000101000: oled_data = 16'b1101110011010110;
				18'b001100100010101000: oled_data = 16'b1101110010010101;
				18'b001100100100101000: oled_data = 16'b1011001101110000;
				18'b001100100110101000: oled_data = 16'b1011001101110001;
				18'b001100101000101000: oled_data = 16'b1100010010110100;
				18'b001100101010101000: oled_data = 16'b1010010100010011;
				18'b001100101100101000: oled_data = 16'b0101101010001001;
				18'b001100101110101000: oled_data = 16'b0100000111000111;
				18'b001100110000101000: oled_data = 16'b0011000101000101;
				18'b001100110010101000: oled_data = 16'b0011000100100101;
				18'b001100110100101000: oled_data = 16'b0100000110100110;
				18'b001100110110101000: oled_data = 16'b0110001011001010;
				18'b001100111000101000: oled_data = 16'b1101011010011001;
				18'b001100111010101000: oled_data = 16'b1110111100111011;
				18'b001100111100101000: oled_data = 16'b1110111100011011;
				18'b001100111110101000: oled_data = 16'b1101010110010111;
				18'b001101000000101000: oled_data = 16'b1100010001010011;
				18'b001101000010101000: oled_data = 16'b1101110011010101;
				18'b001101000100101000: oled_data = 16'b1110010011010110;
				18'b001101000110101000: oled_data = 16'b1100010000110010;
				18'b001101001000101000: oled_data = 16'b0110101010001010;
				18'b001101001010101000: oled_data = 16'b0011100110000110;
				18'b001101001100101000: oled_data = 16'b0011000101000101;
				18'b001101001110101000: oled_data = 16'b0101001000101000;
				18'b001101010000101000: oled_data = 16'b0111001100101101;
				18'b001101010010101000: oled_data = 16'b1010110100010011;
				18'b001101010100101000: oled_data = 16'b1100111000010111;
				18'b001101010110101000: oled_data = 16'b1110011010111010;
				18'b001101011000101000: oled_data = 16'b1110111100111011;
				18'b001101011010101000: oled_data = 16'b1110111101011011;
				18'b001101011100101000: oled_data = 16'b1110111100011011;
				18'b001101011110101000: oled_data = 16'b1110111100011010;
				18'b001101100000101000: oled_data = 16'b1110111100011011;
				18'b001101100010101000: oled_data = 16'b1110111100011010;
				18'b001101100100101000: oled_data = 16'b1110111100011010;
				18'b001101100110101000: oled_data = 16'b1110111100011010;
				18'b001101101000101000: oled_data = 16'b1110111100111011;
				18'b001101101010101000: oled_data = 16'b1100110101110110;
				18'b001101101100101000: oled_data = 16'b1100110000110010;
				18'b001101101110101000: oled_data = 16'b1101110011010101;
				18'b001101110000101000: oled_data = 16'b1101010010010100;
				18'b001101110010101000: oled_data = 16'b1101010001110100;
				18'b001101110100101000: oled_data = 16'b1101010001010100;
				18'b001101110110101000: oled_data = 16'b1101110010110101;
				18'b001101111000101000: oled_data = 16'b1101110011010110;
				18'b001101111010101000: oled_data = 16'b1101110010010101;
				18'b001101111100101000: oled_data = 16'b1101110011110100;
				18'b001101111110101000: oled_data = 16'b1100101111001111;
				18'b001110000000101000: oled_data = 16'b1010101000001000;
				18'b001110000010101000: oled_data = 16'b1011101011101100;
				18'b001110000100101000: oled_data = 16'b1110110011110100;
				18'b001110000110101000: oled_data = 16'b1100101101101110;
				18'b001110001000101000: oled_data = 16'b1011001000101001;
				18'b001110001010101000: oled_data = 16'b1011001001001001;
				18'b001110001100101000: oled_data = 16'b1011001001001001;
				18'b001110001110101000: oled_data = 16'b1011001001001001;
				18'b001110010000101000: oled_data = 16'b1011001001001001;
				18'b001110010010101000: oled_data = 16'b1011001001101010;
				18'b001110010100101000: oled_data = 16'b1100010111111000;
				18'b001110010110101000: oled_data = 16'b1011111100011100;
				18'b001110011000101000: oled_data = 16'b1011111100011100;
				18'b001110011010101000: oled_data = 16'b1011001111101111;
				18'b001110011100101000: oled_data = 16'b1011001000001000;
				18'b001110011110101000: oled_data = 16'b1010101000001000;
				18'b001110100000101000: oled_data = 16'b1010001000001000;
				18'b001110100010101000: oled_data = 16'b1010001000001000;
				18'b001110100100101000: oled_data = 16'b1010101000001000;
				18'b001110100110101000: oled_data = 16'b1010101000001000;
				18'b001100011000101001: oled_data = 16'b1001101111101110;
				18'b001100011010101001: oled_data = 16'b1101110010110101;
				18'b001100011100101001: oled_data = 16'b1101110011010101;
				18'b001100011110101001: oled_data = 16'b1101110011010101;
				18'b001100100000101001: oled_data = 16'b1101110011010101;
				18'b001100100010101001: oled_data = 16'b1101110011010101;
				18'b001100100100101001: oled_data = 16'b1011101111010001;
				18'b001100100110101001: oled_data = 16'b1011001101110001;
				18'b001100101000101001: oled_data = 16'b1100110100010101;
				18'b001100101010101001: oled_data = 16'b1001110010010001;
				18'b001100101100101001: oled_data = 16'b0111001101101101;
				18'b001100101110101001: oled_data = 16'b1000001111101111;
				18'b001100110000101001: oled_data = 16'b1010010011110010;
				18'b001100110010101001: oled_data = 16'b1011110110110110;
				18'b001100110100101001: oled_data = 16'b1101011001011000;
				18'b001100110110101001: oled_data = 16'b1110011011111010;
				18'b001100111000101001: oled_data = 16'b1110011100011010;
				18'b001100111010101001: oled_data = 16'b1110011100011010;
				18'b001100111100101001: oled_data = 16'b1110111100011010;
				18'b001100111110101001: oled_data = 16'b1110111100011011;
				18'b001101000000101001: oled_data = 16'b1101010110110110;
				18'b001101000010101001: oled_data = 16'b1100010010010011;
				18'b001101000100101001: oled_data = 16'b1101110011010101;
				18'b001101000110101001: oled_data = 16'b1101010100010101;
				18'b001101001000101001: oled_data = 16'b1110011010011010;
				18'b001101001010101001: oled_data = 16'b1100010111010110;
				18'b001101001100101001: oled_data = 16'b1000101111101111;
				18'b001101001110101001: oled_data = 16'b0101101001101001;
				18'b001101010000101001: oled_data = 16'b0011100110000110;
				18'b001101010010101001: oled_data = 16'b0011000100100100;
				18'b001101010100101001: oled_data = 16'b0011100101100101;
				18'b001101010110101001: oled_data = 16'b0100101000000111;
				18'b001101011000101001: oled_data = 16'b0110101011101011;
				18'b001101011010101001: oled_data = 16'b1000110000101111;
				18'b001101011100101001: oled_data = 16'b1101011001111000;
				18'b001101011110101001: oled_data = 16'b1110111100011011;
				18'b001101100000101001: oled_data = 16'b1110111100011010;
				18'b001101100010101001: oled_data = 16'b1110111100011010;
				18'b001101100100101001: oled_data = 16'b1110111100011010;
				18'b001101100110101001: oled_data = 16'b1110111100011010;
				18'b001101101000101001: oled_data = 16'b1110111100011010;
				18'b001101101010101001: oled_data = 16'b1111011100011011;
				18'b001101101100101001: oled_data = 16'b1011110010010011;
				18'b001101101110101001: oled_data = 16'b1100010000110010;
				18'b001101110000101001: oled_data = 16'b1101110011110101;
				18'b001101110010101001: oled_data = 16'b1101110011010110;
				18'b001101110100101001: oled_data = 16'b1101110010010101;
				18'b001101110110101001: oled_data = 16'b1101010001110100;
				18'b001101111000101001: oled_data = 16'b1101110010110101;
				18'b001101111010101001: oled_data = 16'b1101110010110101;
				18'b001101111100101001: oled_data = 16'b1101110011110100;
				18'b001101111110101001: oled_data = 16'b1100101110001110;
				18'b001110000000101001: oled_data = 16'b1011001000001000;
				18'b001110000010101001: oled_data = 16'b1100101110101110;
				18'b001110000100101001: oled_data = 16'b1110010011010010;
				18'b001110000110101001: oled_data = 16'b1011101010001010;
				18'b001110001000101001: oled_data = 16'b1011001001001001;
				18'b001110001010101001: oled_data = 16'b1011001001001001;
				18'b001110001100101001: oled_data = 16'b1011001001001001;
				18'b001110001110101001: oled_data = 16'b1011001001001001;
				18'b001110010000101001: oled_data = 16'b1011001000101001;
				18'b001110010010101001: oled_data = 16'b1011001111110000;
				18'b001110010100101001: oled_data = 16'b1100011011111011;
				18'b001110010110101001: oled_data = 16'b1011111011111011;
				18'b001110011000101001: oled_data = 16'b1011111100011100;
				18'b001110011010101001: oled_data = 16'b1011110110110110;
				18'b001110011100101001: oled_data = 16'b1011001001001001;
				18'b001110011110101001: oled_data = 16'b1011001000101000;
				18'b001110100000101001: oled_data = 16'b1011001000101000;
				18'b001110100010101001: oled_data = 16'b1010101000101000;
				18'b001110100100101001: oled_data = 16'b1010101000001000;
				18'b001110100110101001: oled_data = 16'b1010101000001000;
				18'b001100011000101010: oled_data = 16'b1010010000010000;
				18'b001100011010101010: oled_data = 16'b1101110011010101;
				18'b001100011100101010: oled_data = 16'b1101110011010101;
				18'b001100011110101010: oled_data = 16'b1101110011010101;
				18'b001100100000101010: oled_data = 16'b1101110011010101;
				18'b001100100010101010: oled_data = 16'b1101110010110101;
				18'b001100100100101010: oled_data = 16'b1011101110010001;
				18'b001100100110101010: oled_data = 16'b1011001101110001;
				18'b001100101000101010: oled_data = 16'b1101010110010111;
				18'b001100101010101010: oled_data = 16'b1110111100111011;
				18'b001100101100101010: oled_data = 16'b1110111100111011;
				18'b001100101110101010: oled_data = 16'b1110111100111011;
				18'b001100110000101010: oled_data = 16'b1110111100111011;
				18'b001100110010101010: oled_data = 16'b1110111100111011;
				18'b001100110100101010: oled_data = 16'b1110111100011010;
				18'b001100110110101010: oled_data = 16'b1110011100011010;
				18'b001100111000101010: oled_data = 16'b1110011100011010;
				18'b001100111010101010: oled_data = 16'b1110011100011010;
				18'b001100111100101010: oled_data = 16'b1110011100011010;
				18'b001100111110101010: oled_data = 16'b1110011100011010;
				18'b001101000000101010: oled_data = 16'b1110111100011010;
				18'b001101000010101010: oled_data = 16'b1101111000011000;
				18'b001101000100101010: oled_data = 16'b1100110011010100;
				18'b001101000110101010: oled_data = 16'b1101010100010101;
				18'b001101001000101010: oled_data = 16'b1110111011111010;
				18'b001101001010101010: oled_data = 16'b1110111100111011;
				18'b001101001100101010: oled_data = 16'b1110111100111011;
				18'b001101001110101010: oled_data = 16'b1110011011111010;
				18'b001101010000101010: oled_data = 16'b1100111000111000;
				18'b001101010010101010: oled_data = 16'b1010110100110100;
				18'b001101010100101010: oled_data = 16'b1001010001010000;
				18'b001101010110101010: oled_data = 16'b0111001101001100;
				18'b001101011000101010: oled_data = 16'b0101101010101010;
				18'b001101011010101010: oled_data = 16'b0101001001001000;
				18'b001101011100101010: oled_data = 16'b1011110110010101;
				18'b001101011110101010: oled_data = 16'b1110111100111011;
				18'b001101100000101010: oled_data = 16'b1110111100011010;
				18'b001101100010101010: oled_data = 16'b1110111100011010;
				18'b001101100100101010: oled_data = 16'b1110111100011010;
				18'b001101100110101010: oled_data = 16'b1110111100011010;
				18'b001101101000101010: oled_data = 16'b1110111100111011;
				18'b001101101010101010: oled_data = 16'b1101111000110111;
				18'b001101101100101010: oled_data = 16'b1101010100110101;
				18'b001101101110101010: oled_data = 16'b1100110010110011;
				18'b001101110000101010: oled_data = 16'b1101010011010100;
				18'b001101110010101010: oled_data = 16'b1101110011010101;
				18'b001101110100101010: oled_data = 16'b1110010010110101;
				18'b001101110110101010: oled_data = 16'b1101110011010101;
				18'b001101111000101010: oled_data = 16'b1101010001110100;
				18'b001101111010101010: oled_data = 16'b1100110001010100;
				18'b001101111100101010: oled_data = 16'b1101110011010100;
				18'b001101111110101010: oled_data = 16'b1100001101001101;
				18'b001110000000101010: oled_data = 16'b1010101000101000;
				18'b001110000010101010: oled_data = 16'b1101010000110000;
				18'b001110000100101010: oled_data = 16'b1101110000010000;
				18'b001110000110101010: oled_data = 16'b1011001001001001;
				18'b001110001000101010: oled_data = 16'b1011101001001001;
				18'b001110001010101010: oled_data = 16'b1011001001001001;
				18'b001110001100101010: oled_data = 16'b1011001001001001;
				18'b001110001110101010: oled_data = 16'b1011001001001001;
				18'b001110010000101010: oled_data = 16'b1011001001101010;
				18'b001110010010101010: oled_data = 16'b1011110111010111;
				18'b001110010100101010: oled_data = 16'b1011111100011100;
				18'b001110010110101010: oled_data = 16'b1011111011111011;
				18'b001110011000101010: oled_data = 16'b1011111011111100;
				18'b001110011010101010: oled_data = 16'b1100011011011011;
				18'b001110011100101010: oled_data = 16'b1011001101001101;
				18'b001110011110101010: oled_data = 16'b1011001000001000;
				18'b001110100000101010: oled_data = 16'b1011001000101000;
				18'b001110100010101010: oled_data = 16'b1010101000101000;
				18'b001110100100101010: oled_data = 16'b1010101000001000;
				18'b001110100110101010: oled_data = 16'b1010101000001000;
				18'b001100011000101011: oled_data = 16'b1010110000110001;
				18'b001100011010101011: oled_data = 16'b1101110011010101;
				18'b001100011100101011: oled_data = 16'b1101110010110101;
				18'b001100011110101011: oled_data = 16'b1101110010110101;
				18'b001100100000101011: oled_data = 16'b1101110011010101;
				18'b001100100010101011: oled_data = 16'b1101010010010101;
				18'b001100100100101011: oled_data = 16'b1011001101110001;
				18'b001100100110101011: oled_data = 16'b1011001101110001;
				18'b001100101000101011: oled_data = 16'b1101111000111000;
				18'b001100101010101011: oled_data = 16'b1110111100111011;
				18'b001100101100101011: oled_data = 16'b1110011100011010;
				18'b001100101110101011: oled_data = 16'b1110011011111010;
				18'b001100110000101011: oled_data = 16'b1110011100011010;
				18'b001100110010101011: oled_data = 16'b1110111100011010;
				18'b001100110100101011: oled_data = 16'b1110011100011010;
				18'b001100110110101011: oled_data = 16'b1110011011111010;
				18'b001100111000101011: oled_data = 16'b1110011100011010;
				18'b001100111010101011: oled_data = 16'b1110011100011010;
				18'b001100111100101011: oled_data = 16'b1110111100011010;
				18'b001100111110101011: oled_data = 16'b1110111100011010;
				18'b001101000000101011: oled_data = 16'b1110011100011010;
				18'b001101000010101011: oled_data = 16'b1110111100011011;
				18'b001101000100101011: oled_data = 16'b1110011010011010;
				18'b001101000110101011: oled_data = 16'b1101010110110111;
				18'b001101001000101011: oled_data = 16'b1110111100011011;
				18'b001101001010101011: oled_data = 16'b1110011100011010;
				18'b001101001100101011: oled_data = 16'b1110011100011010;
				18'b001101001110101011: oled_data = 16'b1110011100011010;
				18'b001101010000101011: oled_data = 16'b1110111100011010;
				18'b001101010010101011: oled_data = 16'b1110111100011011;
				18'b001101010100101011: oled_data = 16'b1110111100111100;
				18'b001101010110101011: oled_data = 16'b1110111100111011;
				18'b001101011000101011: oled_data = 16'b1110011011111011;
				18'b001101011010101011: oled_data = 16'b1110011011011010;
				18'b001101011100101011: oled_data = 16'b1110011011111010;
				18'b001101011110101011: oled_data = 16'b1110111100011010;
				18'b001101100000101011: oled_data = 16'b1110111100011010;
				18'b001101100010101011: oled_data = 16'b1110111100011010;
				18'b001101100100101011: oled_data = 16'b1110111100011010;
				18'b001101100110101011: oled_data = 16'b1110111100111010;
				18'b001101101000101011: oled_data = 16'b1101111001011000;
				18'b001101101010101011: oled_data = 16'b1101010100110101;
				18'b001101101100101011: oled_data = 16'b1110010101010101;
				18'b001101101110101011: oled_data = 16'b1110010101010110;
				18'b001101110000101011: oled_data = 16'b1101010011110100;
				18'b001101110010101011: oled_data = 16'b1101010011010100;
				18'b001101110100101011: oled_data = 16'b1101010011010101;
				18'b001101110110101011: oled_data = 16'b1101110011010101;
				18'b001101111000101011: oled_data = 16'b1110010011110110;
				18'b001101111010101011: oled_data = 16'b1101110010110101;
				18'b001101111100101011: oled_data = 16'b1101010010110011;
				18'b001101111110101011: oled_data = 16'b1011101100101101;
				18'b001110000000101011: oled_data = 16'b1010101000101001;
				18'b001110000010101011: oled_data = 16'b1101110001110001;
				18'b001110000100101011: oled_data = 16'b1100101101101110;
				18'b001110000110101011: oled_data = 16'b1011001000101001;
				18'b001110001000101011: oled_data = 16'b1011101001001001;
				18'b001110001010101011: oled_data = 16'b1011001001001001;
				18'b001110001100101011: oled_data = 16'b1011001001001001;
				18'b001110001110101011: oled_data = 16'b1011001000101001;
				18'b001110010000101011: oled_data = 16'b1011001101001101;
				18'b001110010010101011: oled_data = 16'b1100011011011011;
				18'b001110010100101011: oled_data = 16'b1011111011111100;
				18'b001110010110101011: oled_data = 16'b1011111011111011;
				18'b001110011000101011: oled_data = 16'b1011111011111100;
				18'b001110011010101011: oled_data = 16'b1100011100111101;
				18'b001110011100101011: oled_data = 16'b1011110100010100;
				18'b001110011110101011: oled_data = 16'b1010101000101001;
				18'b001110100000101011: oled_data = 16'b1011001000101001;
				18'b001110100010101011: oled_data = 16'b1010101000001000;
				18'b001110100100101011: oled_data = 16'b1010101000001000;
				18'b001110100110101011: oled_data = 16'b1010101000001000;
				18'b001100011000101100: oled_data = 16'b1011110001010010;
				18'b001100011010101100: oled_data = 16'b1101110011010101;
				18'b001100011100101100: oled_data = 16'b1101110010110101;
				18'b001100011110101100: oled_data = 16'b1101110010110101;
				18'b001100100000101100: oled_data = 16'b1101110011010110;
				18'b001100100010101100: oled_data = 16'b1100110000110011;
				18'b001100100100101100: oled_data = 16'b1011001101110001;
				18'b001100100110101100: oled_data = 16'b1011001101110000;
				18'b001100101000101100: oled_data = 16'b1101010111110111;
				18'b001100101010101100: oled_data = 16'b1110111100111011;
				18'b001100101100101100: oled_data = 16'b1110011011111010;
				18'b001100101110101100: oled_data = 16'b1110011011111010;
				18'b001100110000101100: oled_data = 16'b1110011011111010;
				18'b001100110010101100: oled_data = 16'b1110011100011010;
				18'b001100110100101100: oled_data = 16'b1110011011111010;
				18'b001100110110101100: oled_data = 16'b1110011011111010;
				18'b001100111000101100: oled_data = 16'b1110111011111010;
				18'b001100111010101100: oled_data = 16'b1110111100011010;
				18'b001100111100101100: oled_data = 16'b1110011100011010;
				18'b001100111110101100: oled_data = 16'b1110011100011010;
				18'b001101000000101100: oled_data = 16'b1110011100011010;
				18'b001101000010101100: oled_data = 16'b1110011011111010;
				18'b001101000100101100: oled_data = 16'b1110111011111011;
				18'b001101000110101100: oled_data = 16'b1110011011111011;
				18'b001101001000101100: oled_data = 16'b1110011011111011;
				18'b001101001010101100: oled_data = 16'b1110011011111011;
				18'b001101001100101100: oled_data = 16'b1110011100011010;
				18'b001101001110101100: oled_data = 16'b1110011100011010;
				18'b001101010000101100: oled_data = 16'b1110011100011010;
				18'b001101010010101100: oled_data = 16'b1110111100011010;
				18'b001101010100101100: oled_data = 16'b1110111100011010;
				18'b001101010110101100: oled_data = 16'b1110111100011010;
				18'b001101011000101100: oled_data = 16'b1110111100011010;
				18'b001101011010101100: oled_data = 16'b1110111100011011;
				18'b001101011100101100: oled_data = 16'b1110111100011011;
				18'b001101011110101100: oled_data = 16'b1110111100011010;
				18'b001101100000101100: oled_data = 16'b1110111100011010;
				18'b001101100010101100: oled_data = 16'b1110111100011010;
				18'b001101100100101100: oled_data = 16'b1110111100011010;
				18'b001101100110101100: oled_data = 16'b1101111000010111;
				18'b001101101000101100: oled_data = 16'b1101010100110100;
				18'b001101101010101100: oled_data = 16'b1101110101010101;
				18'b001101101100101100: oled_data = 16'b1101110101010101;
				18'b001101101110101100: oled_data = 16'b1101110101010101;
				18'b001101110000101100: oled_data = 16'b1101010101110101;
				18'b001101110010101100: oled_data = 16'b1110011011011010;
				18'b001101110100101100: oled_data = 16'b1101111000111000;
				18'b001101110110101100: oled_data = 16'b1100010100110100;
				18'b001101111000101100: oled_data = 16'b1101010100010101;
				18'b001101111010101100: oled_data = 16'b1101110011110101;
				18'b001101111100101100: oled_data = 16'b1101010010110011;
				18'b001101111110101100: oled_data = 16'b1011101100001100;
				18'b001110000000101100: oled_data = 16'b1011001001001010;
				18'b001110000010101100: oled_data = 16'b1101110010010010;
				18'b001110000100101100: oled_data = 16'b1100001011101100;
				18'b001110000110101100: oled_data = 16'b1011001000101001;
				18'b001110001000101100: oled_data = 16'b1011001001001001;
				18'b001110001010101100: oled_data = 16'b1011001001001001;
				18'b001110001100101100: oled_data = 16'b1011001001001001;
				18'b001110001110101100: oled_data = 16'b1011001000101001;
				18'b001110010000101100: oled_data = 16'b1011110010010011;
				18'b001110010010101100: oled_data = 16'b1011111100011100;
				18'b001110010100101100: oled_data = 16'b1011111011111011;
				18'b001110010110101100: oled_data = 16'b1011111011111011;
				18'b001110011000101100: oled_data = 16'b1011111011111100;
				18'b001110011010101100: oled_data = 16'b1100111100111101;
				18'b001110011100101100: oled_data = 16'b1011111001111001;
				18'b001110011110101100: oled_data = 16'b1010101010101011;
				18'b001110100000101100: oled_data = 16'b1010101000101000;
				18'b001110100010101100: oled_data = 16'b1010101000001000;
				18'b001110100100101100: oled_data = 16'b1010101000001000;
				18'b001110100110101100: oled_data = 16'b1010101000001000;
				18'b001100011000101101: oled_data = 16'b1011110001010010;
				18'b001100011010101101: oled_data = 16'b1101110011010101;
				18'b001100011100101101: oled_data = 16'b1101110010110101;
				18'b001100011110101101: oled_data = 16'b1101110010110101;
				18'b001100100000101101: oled_data = 16'b1101110010110110;
				18'b001100100010101101: oled_data = 16'b1100010000010011;
				18'b001100100100101101: oled_data = 16'b1011001101110001;
				18'b001100100110101101: oled_data = 16'b1011001101110001;
				18'b001100101000101101: oled_data = 16'b1011010000110010;
				18'b001100101010101101: oled_data = 16'b1110011011011010;
				18'b001100101100101101: oled_data = 16'b1110111100011010;
				18'b001100101110101101: oled_data = 16'b1110011011111010;
				18'b001100110000101101: oled_data = 16'b1110011011111010;
				18'b001100110010101101: oled_data = 16'b1110011011111010;
				18'b001100110100101101: oled_data = 16'b1110011011111010;
				18'b001100110110101101: oled_data = 16'b1110011011111010;
				18'b001100111000101101: oled_data = 16'b1110011011111010;
				18'b001100111010101101: oled_data = 16'b1110011011111010;
				18'b001100111100101101: oled_data = 16'b1110011011111010;
				18'b001100111110101101: oled_data = 16'b1110011011111010;
				18'b001101000000101101: oled_data = 16'b1110011011111010;
				18'b001101000010101101: oled_data = 16'b1110011011111010;
				18'b001101000100101101: oled_data = 16'b1110011011111010;
				18'b001101000110101101: oled_data = 16'b1110011011111010;
				18'b001101001000101101: oled_data = 16'b1110011011111010;
				18'b001101001010101101: oled_data = 16'b1110011011111010;
				18'b001101001100101101: oled_data = 16'b1110111100011010;
				18'b001101001110101101: oled_data = 16'b1110111100011010;
				18'b001101010000101101: oled_data = 16'b1110111100011010;
				18'b001101010010101101: oled_data = 16'b1110111100011010;
				18'b001101010100101101: oled_data = 16'b1110111100011010;
				18'b001101010110101101: oled_data = 16'b1110111100011010;
				18'b001101011000101101: oled_data = 16'b1110111100011010;
				18'b001101011010101101: oled_data = 16'b1110111100011010;
				18'b001101011100101101: oled_data = 16'b1110111100011010;
				18'b001101011110101101: oled_data = 16'b1110111100011010;
				18'b001101100000101101: oled_data = 16'b1110111100111010;
				18'b001101100010101101: oled_data = 16'b1110111100011010;
				18'b001101100100101101: oled_data = 16'b1101010111010110;
				18'b001101100110101101: oled_data = 16'b1101010100010100;
				18'b001101101000101101: oled_data = 16'b1101110100010101;
				18'b001101101010101101: oled_data = 16'b1101110100110101;
				18'b001101101100101101: oled_data = 16'b1110010101010101;
				18'b001101101110101101: oled_data = 16'b1101010101010101;
				18'b001101110000101101: oled_data = 16'b1101111001011000;
				18'b001101110010101101: oled_data = 16'b1110111011111010;
				18'b001101110100101101: oled_data = 16'b1110011010111001;
				18'b001101110110101101: oled_data = 16'b1110011010111001;
				18'b001101111000101101: oled_data = 16'b1110011010011001;
				18'b001101111010101101: oled_data = 16'b1101010111010111;
				18'b001101111100101101: oled_data = 16'b1100110100010100;
				18'b001101111110101101: oled_data = 16'b1011101011101100;
				18'b001110000000101101: oled_data = 16'b1011001001001010;
				18'b001110000010101101: oled_data = 16'b1101110001110001;
				18'b001110000100101101: oled_data = 16'b1011101010001011;
				18'b001110000110101101: oled_data = 16'b1011001001001001;
				18'b001110001000101101: oled_data = 16'b1011001001001001;
				18'b001110001010101101: oled_data = 16'b1011001001001001;
				18'b001110001100101101: oled_data = 16'b1011001000101001;
				18'b001110001110101101: oled_data = 16'b1011001001001001;
				18'b001110010000101101: oled_data = 16'b1100010111010111;
				18'b001110010010101101: oled_data = 16'b1011111100011100;
				18'b001110010100101101: oled_data = 16'b1011111011111011;
				18'b001110010110101101: oled_data = 16'b1011111011111011;
				18'b001110011000101101: oled_data = 16'b1011111011111011;
				18'b001110011010101101: oled_data = 16'b1100111100011100;
				18'b001110011100101101: oled_data = 16'b1011111011111011;
				18'b001110011110101101: oled_data = 16'b1011001110101110;
				18'b001110100000101101: oled_data = 16'b1010101000001000;
				18'b001110100010101101: oled_data = 16'b1010101000001000;
				18'b001110100100101101: oled_data = 16'b1010101000001000;
				18'b001110100110101101: oled_data = 16'b1010101000001000;
				18'b001100011000101110: oled_data = 16'b1011010000010001;
				18'b001100011010101110: oled_data = 16'b1101110010110101;
				18'b001100011100101110: oled_data = 16'b1101110010110101;
				18'b001100011110101110: oled_data = 16'b1101110010110101;
				18'b001100100000101110: oled_data = 16'b1101110010110101;
				18'b001100100010101110: oled_data = 16'b1100001111110010;
				18'b001100100100101110: oled_data = 16'b1011001101110001;
				18'b001100100110101110: oled_data = 16'b1011001110010001;
				18'b001100101000101110: oled_data = 16'b1010101101010000;
				18'b001100101010101110: oled_data = 16'b1011010001010010;
				18'b001100101100101110: oled_data = 16'b1110011010111010;
				18'b001100101110101110: oled_data = 16'b1110011100011010;
				18'b001100110000101110: oled_data = 16'b1110011011111010;
				18'b001100110010101110: oled_data = 16'b1110011100011010;
				18'b001100110100101110: oled_data = 16'b1110011100011010;
				18'b001100110110101110: oled_data = 16'b1110011011111010;
				18'b001100111000101110: oled_data = 16'b1110011011111010;
				18'b001100111010101110: oled_data = 16'b1110011011111010;
				18'b001100111100101110: oled_data = 16'b1110011011111010;
				18'b001100111110101110: oled_data = 16'b1110011011111010;
				18'b001101000000101110: oled_data = 16'b1110011011111010;
				18'b001101000010101110: oled_data = 16'b1110011011111010;
				18'b001101000100101110: oled_data = 16'b1110011011111010;
				18'b001101000110101110: oled_data = 16'b1110011011111010;
				18'b001101001000101110: oled_data = 16'b1110011011111010;
				18'b001101001010101110: oled_data = 16'b1110011011111010;
				18'b001101001100101110: oled_data = 16'b1110011100011010;
				18'b001101001110101110: oled_data = 16'b1110011100011010;
				18'b001101010000101110: oled_data = 16'b1110011100011010;
				18'b001101010010101110: oled_data = 16'b1110011100011010;
				18'b001101010100101110: oled_data = 16'b1110011100011010;
				18'b001101010110101110: oled_data = 16'b1110111100011010;
				18'b001101011000101110: oled_data = 16'b1110111100011010;
				18'b001101011010101110: oled_data = 16'b1110111100011010;
				18'b001101011100101110: oled_data = 16'b1110011100011010;
				18'b001101011110101110: oled_data = 16'b1110111100011010;
				18'b001101100000101110: oled_data = 16'b1110011010111001;
				18'b001101100010101110: oled_data = 16'b1100010100010011;
				18'b001101100100101110: oled_data = 16'b1101010011110100;
				18'b001101100110101110: oled_data = 16'b1101010011110100;
				18'b001101101000101110: oled_data = 16'b1101010011110101;
				18'b001101101010101110: oled_data = 16'b1101110100110101;
				18'b001101101100101110: oled_data = 16'b1101110100110101;
				18'b001101101110101110: oled_data = 16'b1101010111010111;
				18'b001101110000101110: oled_data = 16'b1110111011111010;
				18'b001101110010101110: oled_data = 16'b1110011011011001;
				18'b001101110100101110: oled_data = 16'b1101111010011000;
				18'b001101110110101110: oled_data = 16'b1110111011111010;
				18'b001101111000101110: oled_data = 16'b1110011100011010;
				18'b001101111010101110: oled_data = 16'b1110111100011011;
				18'b001101111100101110: oled_data = 16'b1101111000110111;
				18'b001101111110101110: oled_data = 16'b1011001011001011;
				18'b001110000000101110: oled_data = 16'b1011001001101010;
				18'b001110000010101110: oled_data = 16'b1101010000110000;
				18'b001110000100101110: oled_data = 16'b1011101001101010;
				18'b001110000110101110: oled_data = 16'b1011001001001001;
				18'b001110001000101110: oled_data = 16'b1011001001001001;
				18'b001110001010101110: oled_data = 16'b1011001001001001;
				18'b001110001100101110: oled_data = 16'b1011001000101001;
				18'b001110001110101110: oled_data = 16'b1011001010101011;
				18'b001110010000101110: oled_data = 16'b1100011001111010;
				18'b001110010010101110: oled_data = 16'b1011111011111100;
				18'b001110010100101110: oled_data = 16'b1011111011011011;
				18'b001110010110101110: oled_data = 16'b1011111011111011;
				18'b001110011000101110: oled_data = 16'b1011111011111011;
				18'b001110011010101110: oled_data = 16'b1100111100011100;
				18'b001110011100101110: oled_data = 16'b1011111100011100;
				18'b001110011110101110: oled_data = 16'b1011010010110010;
				18'b001110100000101110: oled_data = 16'b1010100111101000;
				18'b001110100010101110: oled_data = 16'b1010101000001000;
				18'b001110100100101110: oled_data = 16'b1010101000001000;
				18'b001110100110101110: oled_data = 16'b1010101000001000;
				18'b001100011000101111: oled_data = 16'b1010101111110001;
				18'b001100011010101111: oled_data = 16'b1101110010010101;
				18'b001100011100101111: oled_data = 16'b1101010001110100;
				18'b001100011110101111: oled_data = 16'b1101010010010100;
				18'b001100100000101111: oled_data = 16'b1101110010110101;
				18'b001100100010101111: oled_data = 16'b1100001111010010;
				18'b001100100100101111: oled_data = 16'b1011001101010000;
				18'b001100100110101111: oled_data = 16'b1011001101110000;
				18'b001100101000101111: oled_data = 16'b1010101100110000;
				18'b001100101010101111: oled_data = 16'b1010101100110000;
				18'b001100101100101111: oled_data = 16'b1011010000010010;
				18'b001100101110101111: oled_data = 16'b1110011001111001;
				18'b001100110000101111: oled_data = 16'b1110111100011010;
				18'b001100110010101111: oled_data = 16'b1110011100011010;
				18'b001100110100101111: oled_data = 16'b1110011011111010;
				18'b001100110110101111: oled_data = 16'b1110011011111010;
				18'b001100111000101111: oled_data = 16'b1110011011111010;
				18'b001100111010101111: oled_data = 16'b1110011011111010;
				18'b001100111100101111: oled_data = 16'b1110011011111010;
				18'b001100111110101111: oled_data = 16'b1110011011111010;
				18'b001101000000101111: oled_data = 16'b1110011011111010;
				18'b001101000010101111: oled_data = 16'b1110011011111010;
				18'b001101000100101111: oled_data = 16'b1110011011111010;
				18'b001101000110101111: oled_data = 16'b1110011011111010;
				18'b001101001000101111: oled_data = 16'b1110011011111010;
				18'b001101001010101111: oled_data = 16'b1110011011111010;
				18'b001101001100101111: oled_data = 16'b1110011011111010;
				18'b001101001110101111: oled_data = 16'b1110011011111010;
				18'b001101010000101111: oled_data = 16'b1110011011111010;
				18'b001101010010101111: oled_data = 16'b1110011100011010;
				18'b001101010100101111: oled_data = 16'b1110011100011010;
				18'b001101010110101111: oled_data = 16'b1110011100011010;
				18'b001101011000101111: oled_data = 16'b1110011100011010;
				18'b001101011010101111: oled_data = 16'b1110011100011010;
				18'b001101011100101111: oled_data = 16'b1110011100011010;
				18'b001101011110101111: oled_data = 16'b1101011000010111;
				18'b001101100000101111: oled_data = 16'b1011010000010000;
				18'b001101100010101111: oled_data = 16'b1100010000010001;
				18'b001101100100101111: oled_data = 16'b1101110100110101;
				18'b001101100110101111: oled_data = 16'b1101010011010100;
				18'b001101101000101111: oled_data = 16'b1101110100010101;
				18'b001101101010101111: oled_data = 16'b1101110100010110;
				18'b001101101100101111: oled_data = 16'b1101010100010101;
				18'b001101101110101111: oled_data = 16'b1101110111110111;
				18'b001101110000101111: oled_data = 16'b1110011011111010;
				18'b001101110010101111: oled_data = 16'b1101111010011000;
				18'b001101110100101111: oled_data = 16'b1110011011111010;
				18'b001101110110101111: oled_data = 16'b1110111011111010;
				18'b001101111000101111: oled_data = 16'b1110011011111010;
				18'b001101111010101111: oled_data = 16'b1110011100011010;
				18'b001101111100101111: oled_data = 16'b1110011011111001;
				18'b001101111110101111: oled_data = 16'b1010101100101100;
				18'b001110000000101111: oled_data = 16'b1011001001101010;
				18'b001110000010101111: oled_data = 16'b1100101111101111;
				18'b001110000100101111: oled_data = 16'b1011001001001001;
				18'b001110000110101111: oled_data = 16'b1011001001001001;
				18'b001110001000101111: oled_data = 16'b1011001001101001;
				18'b001110001010101111: oled_data = 16'b1011001001001001;
				18'b001110001100101111: oled_data = 16'b1011001000101000;
				18'b001110001110101111: oled_data = 16'b1011101011101100;
				18'b001110010000101111: oled_data = 16'b1100011010111011;
				18'b001110010010101111: oled_data = 16'b1011111011011100;
				18'b001110010100101111: oled_data = 16'b1011111011011011;
				18'b001110010110101111: oled_data = 16'b1011111011111100;
				18'b001110011000101111: oled_data = 16'b1011111011111100;
				18'b001110011010101111: oled_data = 16'b1011111011111100;
				18'b001110011100101111: oled_data = 16'b1011111100011100;
				18'b001110011110101111: oled_data = 16'b1011110100010100;
				18'b001110100000101111: oled_data = 16'b1010100111101000;
				18'b001110100010101111: oled_data = 16'b1010100111101000;
				18'b001110100100101111: oled_data = 16'b1010101000001000;
				18'b001110100110101111: oled_data = 16'b1010100111101000;
				18'b001100011000110000: oled_data = 16'b1010101111110001;
				18'b001100011010110000: oled_data = 16'b1101110001110101;
				18'b001100011100110000: oled_data = 16'b1100110001010011;
				18'b001100011110110000: oled_data = 16'b1100110000110011;
				18'b001100100000110000: oled_data = 16'b1101010010010101;
				18'b001100100010110000: oled_data = 16'b1011101110110001;
				18'b001100100100110000: oled_data = 16'b1010101100110000;
				18'b001100100110110000: oled_data = 16'b1011001101010000;
				18'b001100101000110000: oled_data = 16'b1010101100001111;
				18'b001100101010110000: oled_data = 16'b1011001101010000;
				18'b001100101100110000: oled_data = 16'b1010001011101111;
				18'b001100101110110000: oled_data = 16'b1011001101110000;
				18'b001100110000110000: oled_data = 16'b1100110101010110;
				18'b001100110010110000: oled_data = 16'b1110011011111010;
				18'b001100110100110000: oled_data = 16'b1110011011111010;
				18'b001100110110110000: oled_data = 16'b1110011011111010;
				18'b001100111000110000: oled_data = 16'b1110011011011001;
				18'b001100111010110000: oled_data = 16'b1110011011011001;
				18'b001100111100110000: oled_data = 16'b1110011011011001;
				18'b001100111110110000: oled_data = 16'b1110011011011001;
				18'b001101000000110000: oled_data = 16'b1110011011011001;
				18'b001101000010110000: oled_data = 16'b1110011011011001;
				18'b001101000100110000: oled_data = 16'b1110011011011001;
				18'b001101000110110000: oled_data = 16'b1110011011111010;
				18'b001101001000110000: oled_data = 16'b1110011011111010;
				18'b001101001010110000: oled_data = 16'b1110011011111010;
				18'b001101001100110000: oled_data = 16'b1110011011111010;
				18'b001101001110110000: oled_data = 16'b1110011011111010;
				18'b001101010000110000: oled_data = 16'b1110011011111010;
				18'b001101010010110000: oled_data = 16'b1110011011111010;
				18'b001101010100110000: oled_data = 16'b1110011011111010;
				18'b001101010110110000: oled_data = 16'b1110011100011010;
				18'b001101011000110000: oled_data = 16'b1110111100011010;
				18'b001101011010110000: oled_data = 16'b1101111010011000;
				18'b001101011100110000: oled_data = 16'b1100010011110011;
				18'b001101011110110000: oled_data = 16'b1011001110101111;
				18'b001101100000110000: oled_data = 16'b1011101110110000;
				18'b001101100010110000: oled_data = 16'b1101110011010100;
				18'b001101100100110000: oled_data = 16'b1101010010110011;
				18'b001101100110110000: oled_data = 16'b1101110011110100;
				18'b001101101000110000: oled_data = 16'b1101110100010101;
				18'b001101101010110000: oled_data = 16'b1101110100010101;
				18'b001101101100110000: oled_data = 16'b1101110100010101;
				18'b001101101110110000: oled_data = 16'b1100110101010101;
				18'b001101110000110000: oled_data = 16'b1101111000111000;
				18'b001101110010110000: oled_data = 16'b1110011010111001;
				18'b001101110100110000: oled_data = 16'b1110011011111010;
				18'b001101110110110000: oled_data = 16'b1110011011111010;
				18'b001101111000110000: oled_data = 16'b1110011011111010;
				18'b001101111010110000: oled_data = 16'b1110011100011010;
				18'b001101111100110000: oled_data = 16'b1110011011011001;
				18'b001101111110110000: oled_data = 16'b1011001110101110;
				18'b001110000000110000: oled_data = 16'b1011001001101010;
				18'b001110000010110000: oled_data = 16'b1100101110001110;
				18'b001110000100110000: oled_data = 16'b1011001000101001;
				18'b001110000110110000: oled_data = 16'b1011001000101001;
				18'b001110001000110000: oled_data = 16'b1100101101101101;
				18'b001110001010110000: oled_data = 16'b1011101001101010;
				18'b001110001100110000: oled_data = 16'b1011001000101000;
				18'b001110001110110000: oled_data = 16'b1011101100001100;
				18'b001110010000110000: oled_data = 16'b1100011011011011;
				18'b001110010010110000: oled_data = 16'b1011111011111100;
				18'b001110010100110000: oled_data = 16'b1011111011011100;
				18'b001110010110110000: oled_data = 16'b1011011010011010;
				18'b001110011000110000: oled_data = 16'b1010011001011001;
				18'b001110011010110000: oled_data = 16'b1011011010111011;
				18'b001110011100110000: oled_data = 16'b1011111100011100;
				18'b001110011110110000: oled_data = 16'b1011110100010100;
				18'b001110100000110000: oled_data = 16'b1010100111001000;
				18'b001110100010110000: oled_data = 16'b1001100111000111;
				18'b001110100100110000: oled_data = 16'b1001100111000111;
				18'b001110100110110000: oled_data = 16'b1001100111000111;
				18'b001100011000110001: oled_data = 16'b1010001110110000;
				18'b001100011010110001: oled_data = 16'b1101010001110101;
				18'b001100011100110001: oled_data = 16'b1100110001010011;
				18'b001100011110110001: oled_data = 16'b1100010000010010;
				18'b001100100000110001: oled_data = 16'b1101010001110100;
				18'b001100100010110001: oled_data = 16'b1011101110010001;
				18'b001100100100110001: oled_data = 16'b1010101100101111;
				18'b001100100110110001: oled_data = 16'b1010101100101111;
				18'b001100101000110001: oled_data = 16'b1010101100001111;
				18'b001100101010110001: oled_data = 16'b1010101100110000;
				18'b001100101100110001: oled_data = 16'b1010001011001110;
				18'b001100101110110001: oled_data = 16'b1010001011101110;
				18'b001100110000110001: oled_data = 16'b1010001100001111;
				18'b001100110010110001: oled_data = 16'b1011010001010010;
				18'b001100110100110001: oled_data = 16'b1101010110110111;
				18'b001100110110110001: oled_data = 16'b1110011010111010;
				18'b001100111000110001: oled_data = 16'b1110111100011010;
				18'b001100111010110001: oled_data = 16'b1110011011111010;
				18'b001100111100110001: oled_data = 16'b1110011011011010;
				18'b001100111110110001: oled_data = 16'b1110011011011010;
				18'b001101000000110001: oled_data = 16'b1110011011011001;
				18'b001101000010110001: oled_data = 16'b1110011011011010;
				18'b001101000100110001: oled_data = 16'b1110011011011010;
				18'b001101000110110001: oled_data = 16'b1110011011011010;
				18'b001101001000110001: oled_data = 16'b1110011011011010;
				18'b001101001010110001: oled_data = 16'b1110011011011010;
				18'b001101001100110001: oled_data = 16'b1110011011011010;
				18'b001101001110110001: oled_data = 16'b1110011011111010;
				18'b001101010000110001: oled_data = 16'b1110011011111010;
				18'b001101010010110001: oled_data = 16'b1110011100011010;
				18'b001101010100110001: oled_data = 16'b1110011100011010;
				18'b001101010110110001: oled_data = 16'b1101111010011000;
				18'b001101011000110001: oled_data = 16'b1100010100110100;
				18'b001101011010110001: oled_data = 16'b1011001111010000;
				18'b001101011100110001: oled_data = 16'b1011101110001111;
				18'b001101011110110001: oled_data = 16'b1011101110110000;
				18'b001101100000110001: oled_data = 16'b1100110001110010;
				18'b001101100010110001: oled_data = 16'b1101110011110100;
				18'b001101100100110001: oled_data = 16'b1100110010010011;
				18'b001101100110110001: oled_data = 16'b1101110100010101;
				18'b001101101000110001: oled_data = 16'b1101110100010101;
				18'b001101101010110001: oled_data = 16'b1101110100010101;
				18'b001101101100110001: oled_data = 16'b1101110100010101;
				18'b001101101110110001: oled_data = 16'b1101010100110101;
				18'b001101110000110001: oled_data = 16'b1100110100010100;
				18'b001101110010110001: oled_data = 16'b1110011001011000;
				18'b001101110100110001: oled_data = 16'b1110111100011010;
				18'b001101110110110001: oled_data = 16'b1110011011111010;
				18'b001101111000110001: oled_data = 16'b1110011011111010;
				18'b001101111010110001: oled_data = 16'b1110011011111010;
				18'b001101111100110001: oled_data = 16'b1101111001111000;
				18'b001101111110110001: oled_data = 16'b1011001111001110;
				18'b001110000000110001: oled_data = 16'b1011001001001001;
				18'b001110000010110001: oled_data = 16'b1100001101001101;
				18'b001110000100110001: oled_data = 16'b1011001000101001;
				18'b001110000110110001: oled_data = 16'b1011001001001001;
				18'b001110001000110001: oled_data = 16'b1100101101101101;
				18'b001110001010110001: oled_data = 16'b1011001001001001;
				18'b001110001100110001: oled_data = 16'b1011001000001000;
				18'b001110001110110001: oled_data = 16'b1011101011001011;
				18'b001110010000110001: oled_data = 16'b1100011010111010;
				18'b001110010010110001: oled_data = 16'b1011111011111100;
				18'b001110010100110001: oled_data = 16'b1010111010011011;
				18'b001110010110110001: oled_data = 16'b1001010111011000;
				18'b001110011000110001: oled_data = 16'b1001010110110111;
				18'b001110011010110001: oled_data = 16'b1010111001111010;
				18'b001110011100110001: oled_data = 16'b1011011011111100;
				18'b001110011110110001: oled_data = 16'b1011010001110010;
				18'b001110100000110001: oled_data = 16'b1010000110100111;
				18'b001110100010110001: oled_data = 16'b1010100111101000;
				18'b001110100100110001: oled_data = 16'b1010000111101000;
				18'b001110100110110001: oled_data = 16'b1010000111000111;
				18'b001100011000110010: oled_data = 16'b1000001100001101;
				18'b001100011010110010: oled_data = 16'b1101010001110101;
				18'b001100011100110010: oled_data = 16'b1100110000110011;
				18'b001100011110110010: oled_data = 16'b1100001111110010;
				18'b001100100000110010: oled_data = 16'b1100110000110011;
				18'b001100100010110010: oled_data = 16'b1011001110010001;
				18'b001100100100110010: oled_data = 16'b1010101100101111;
				18'b001100100110110010: oled_data = 16'b1010001011001110;
				18'b001100101000110010: oled_data = 16'b1010001011101111;
				18'b001100101010110010: oled_data = 16'b1010101100001111;
				18'b001100101100110010: oled_data = 16'b1001101010101110;
				18'b001100101110110010: oled_data = 16'b1010001011001110;
				18'b001100110000110010: oled_data = 16'b1010101100001111;
				18'b001100110010110010: oled_data = 16'b1010101101001111;
				18'b001100110100110010: oled_data = 16'b1010101101001111;
				18'b001100110110110010: oled_data = 16'b1011001111110001;
				18'b001100111000110010: oled_data = 16'b1100010011110100;
				18'b001100111010110010: oled_data = 16'b1101010111010110;
				18'b001100111100110010: oled_data = 16'b1110011001111001;
				18'b001100111110110010: oled_data = 16'b1110111010111010;
				18'b001101000000110010: oled_data = 16'b1110111011111010;
				18'b001101000010110010: oled_data = 16'b1110111011111010;
				18'b001101000100110010: oled_data = 16'b1110011011111010;
				18'b001101000110110010: oled_data = 16'b1110111011111010;
				18'b001101001000110010: oled_data = 16'b1110011011011010;
				18'b001101001010110010: oled_data = 16'b1110011010111001;
				18'b001101001100110010: oled_data = 16'b1110011010111001;
				18'b001101001110110010: oled_data = 16'b1110011011111010;
				18'b001101010000110010: oled_data = 16'b1101111010111001;
				18'b001101010010110010: oled_data = 16'b1101010111110110;
				18'b001101010100110010: oled_data = 16'b1011110011010011;
				18'b001101010110110010: oled_data = 16'b1010101110101111;
				18'b001101011000110010: oled_data = 16'b1011001110001111;
				18'b001101011010110010: oled_data = 16'b1011101110110000;
				18'b001101011100110010: oled_data = 16'b1011101111010000;
				18'b001101011110110010: oled_data = 16'b1100110001010010;
				18'b001101100000110010: oled_data = 16'b1101010010110011;
				18'b001101100010110010: oled_data = 16'b1100110010010011;
				18'b001101100100110010: oled_data = 16'b1101010011110100;
				18'b001101100110110010: oled_data = 16'b1101110011110101;
				18'b001101101000110010: oled_data = 16'b1101110011110101;
				18'b001101101010110010: oled_data = 16'b1101110011110101;
				18'b001101101100110010: oled_data = 16'b1101110100010101;
				18'b001101101110110010: oled_data = 16'b1101110100010101;
				18'b001101110000110010: oled_data = 16'b1101010011110100;
				18'b001101110010110010: oled_data = 16'b1100110011110100;
				18'b001101110100110010: oled_data = 16'b1100110110010110;
				18'b001101110110110010: oled_data = 16'b1110011011011010;
				18'b001101111000110010: oled_data = 16'b1110111100011010;
				18'b001101111010110010: oled_data = 16'b1110011011011001;
				18'b001101111100110010: oled_data = 16'b1110011011111010;
				18'b001101111110110010: oled_data = 16'b1011001110101110;
				18'b001110000000110010: oled_data = 16'b1011001001001001;
				18'b001110000010110010: oled_data = 16'b1100001100101100;
				18'b001110000100110010: oled_data = 16'b1011001000101001;
				18'b001110000110110010: oled_data = 16'b1011001001001001;
				18'b001110001000110010: oled_data = 16'b1011101010101010;
				18'b001110001010110010: oled_data = 16'b1011001000101000;
				18'b001110001100110010: oled_data = 16'b1011001000001000;
				18'b001110001110110010: oled_data = 16'b1011001001001001;
				18'b001110010000110010: oled_data = 16'b1100011000111000;
				18'b001110010010110010: oled_data = 16'b1011111011111100;
				18'b001110010100110010: oled_data = 16'b1001111000011000;
				18'b001110010110110010: oled_data = 16'b1000110110110111;
				18'b001110011000110010: oled_data = 16'b1000110110110111;
				18'b001110011010110010: oled_data = 16'b1001010110111000;
				18'b001110011100110010: oled_data = 16'b1010111001111010;
				18'b001110011110110010: oled_data = 16'b1010101110001110;
				18'b001110100000110010: oled_data = 16'b1010000110100111;
				18'b001110100010110010: oled_data = 16'b1010000111100111;
				18'b001110100100110010: oled_data = 16'b1010000111000111;
				18'b001110100110110010: oled_data = 16'b1010000111000111;
				18'b001100011000110011: oled_data = 16'b0110101001001010;
				18'b001100011010110011: oled_data = 16'b1100110001010100;
				18'b001100011100110011: oled_data = 16'b1100110000010011;
				18'b001100011110110011: oled_data = 16'b1100001111010010;
				18'b001100100000110011: oled_data = 16'b1100110000010011;
				18'b001100100010110011: oled_data = 16'b1100001111110010;
				18'b001100100100110011: oled_data = 16'b1010101100110000;
				18'b001100100110110011: oled_data = 16'b1001101010101101;
				18'b001100101000110011: oled_data = 16'b1010001011101110;
				18'b001100101010110011: oled_data = 16'b1010001011101111;
				18'b001100101100110011: oled_data = 16'b1001101010001101;
				18'b001100101110110011: oled_data = 16'b1001101010101101;
				18'b001100110000110011: oled_data = 16'b1010101100101111;
				18'b001100110010110011: oled_data = 16'b1010101100101110;
				18'b001100110100110011: oled_data = 16'b1010001100001110;
				18'b001100110110110011: oled_data = 16'b1010101100001110;
				18'b001100111000110011: oled_data = 16'b1010101100001110;
				18'b001100111010110011: oled_data = 16'b1010101100101111;
				18'b001100111100110011: oled_data = 16'b1010101110110000;
				18'b001100111110110011: oled_data = 16'b1011110000010001;
				18'b001101000000110011: oled_data = 16'b1100010011110100;
				18'b001101000010110011: oled_data = 16'b1101010110010101;
				18'b001101000100110011: oled_data = 16'b1101010111010110;
				18'b001101000110110011: oled_data = 16'b1100110111010110;
				18'b001101001000110011: oled_data = 16'b1100111000110111;
				18'b001101001010110011: oled_data = 16'b1101011001111000;
				18'b001101001100110011: oled_data = 16'b1101011001010111;
				18'b001101001110110011: oled_data = 16'b1011010011010010;
				18'b001101010000110011: oled_data = 16'b1010101111001111;
				18'b001101010010110011: oled_data = 16'b1011001101101111;
				18'b001101010100110011: oled_data = 16'b1011001101101111;
				18'b001101010110110011: oled_data = 16'b1011001101101110;
				18'b001101011000110011: oled_data = 16'b1011001101101111;
				18'b001101011010110011: oled_data = 16'b1011001110110000;
				18'b001101011100110011: oled_data = 16'b1100110001010010;
				18'b001101011110110011: oled_data = 16'b1101010010110100;
				18'b001101100000110011: oled_data = 16'b1100010000010001;
				18'b001101100010110011: oled_data = 16'b1101010010110011;
				18'b001101100100110011: oled_data = 16'b1101010011110100;
				18'b001101100110110011: oled_data = 16'b1101010011110100;
				18'b001101101000110011: oled_data = 16'b1101010011110100;
				18'b001101101010110011: oled_data = 16'b1101010011110100;
				18'b001101101100110011: oled_data = 16'b1101010011110101;
				18'b001101101110110011: oled_data = 16'b1101010011110101;
				18'b001101110000110011: oled_data = 16'b1101010011010101;
				18'b001101110010110011: oled_data = 16'b1101010011010100;
				18'b001101110100110011: oled_data = 16'b0110101000101001;
				18'b001101110110110011: oled_data = 16'b0101001000101000;
				18'b001101111000110011: oled_data = 16'b1011010101010011;
				18'b001101111010110011: oled_data = 16'b1110011011011001;
				18'b001101111100110011: oled_data = 16'b1010010011010001;
				18'b001101111110110011: oled_data = 16'b1000001001001000;
				18'b001110000000110011: oled_data = 16'b1011001001001001;
				18'b001110000010110011: oled_data = 16'b1011101100001100;
				18'b001110000100110011: oled_data = 16'b1010101000001000;
				18'b001110000110110011: oled_data = 16'b1011001000001000;
				18'b001110001000110011: oled_data = 16'b1011001000001000;
				18'b001110001010110011: oled_data = 16'b1011001000001000;
				18'b001110001100110011: oled_data = 16'b1010101000001000;
				18'b001110001110110011: oled_data = 16'b1011001000001000;
				18'b001110010000110011: oled_data = 16'b1011110001110001;
				18'b001110010010110011: oled_data = 16'b1011111011111011;
				18'b001110010100110011: oled_data = 16'b1001010111010111;
				18'b001110010110110011: oled_data = 16'b1000110101110110;
				18'b001110011000110011: oled_data = 16'b1000110101110110;
				18'b001110011010110011: oled_data = 16'b1000110110010111;
				18'b001110011100110011: oled_data = 16'b1010010110010110;
				18'b001110011110110011: oled_data = 16'b1001101000101001;
				18'b001110100000110011: oled_data = 16'b1010000111000111;
				18'b001110100010110011: oled_data = 16'b1001100111000111;
				18'b001110100100110011: oled_data = 16'b1001100111000111;
				18'b001110100110110011: oled_data = 16'b1001100111000111;
				18'b001100011000110100: oled_data = 16'b0100100111001000;
				18'b001100011010110100: oled_data = 16'b1011101111110010;
				18'b001100011100110100: oled_data = 16'b1100101111110011;
				18'b001100011110110100: oled_data = 16'b1100001111110010;
				18'b001100100000110100: oled_data = 16'b1011101110110010;
				18'b001100100010110100: oled_data = 16'b1100001111010010;
				18'b001100100100110100: oled_data = 16'b1100001111010010;
				18'b001100100110110100: oled_data = 16'b1010001011001110;
				18'b001100101000110100: oled_data = 16'b1010001011001110;
				18'b001100101010110100: oled_data = 16'b1010001011101111;
				18'b001100101100110100: oled_data = 16'b1001101010001101;
				18'b001100101110110100: oled_data = 16'b1001001010001101;
				18'b001100110000110100: oled_data = 16'b1011001101010000;
				18'b001100110010110100: oled_data = 16'b1011001101101111;
				18'b001100110100110100: oled_data = 16'b1010101100101110;
				18'b001100110110110100: oled_data = 16'b1010101100001110;
				18'b001100111000110100: oled_data = 16'b1010101100101110;
				18'b001100111010110100: oled_data = 16'b1011001110010000;
				18'b001100111100110100: oled_data = 16'b1011001110010000;
				18'b001100111110110100: oled_data = 16'b1011001101110000;
				18'b001101000000110100: oled_data = 16'b1011001101101111;
				18'b001101000010110100: oled_data = 16'b1010101101001110;
				18'b001101000100110100: oled_data = 16'b1010101100101110;
				18'b001101000110110100: oled_data = 16'b1011010001110001;
				18'b001101001000110100: oled_data = 16'b1101011001111000;
				18'b001101001010110100: oled_data = 16'b1101111010111001;
				18'b001101001100110100: oled_data = 16'b1101111010111001;
				18'b001101001110110100: oled_data = 16'b1101011000010111;
				18'b001101010000110100: oled_data = 16'b1011010000110001;
				18'b001101010010110100: oled_data = 16'b1011001101101111;
				18'b001101010100110100: oled_data = 16'b1010101101001110;
				18'b001101010110110100: oled_data = 16'b1010101101001110;
				18'b001101011000110100: oled_data = 16'b1011001110101111;
				18'b001101011010110100: oled_data = 16'b1100010000110001;
				18'b001101011100110100: oled_data = 16'b1100110001010010;
				18'b001101011110110100: oled_data = 16'b1100110001110010;
				18'b001101100000110100: oled_data = 16'b1100010001010001;
				18'b001101100010110100: oled_data = 16'b1101010010110011;
				18'b001101100100110100: oled_data = 16'b1101010011010100;
				18'b001101100110110100: oled_data = 16'b1101010011010100;
				18'b001101101000110100: oled_data = 16'b1101010011010100;
				18'b001101101010110100: oled_data = 16'b1101010011010100;
				18'b001101101100110100: oled_data = 16'b1101010011010100;
				18'b001101101110110100: oled_data = 16'b1101010011010100;
				18'b001101110000110100: oled_data = 16'b1101010011010100;
				18'b001101110010110100: oled_data = 16'b1100010001010010;
				18'b001101110100110100: oled_data = 16'b0011000011100011;
				18'b001101110110110100: oled_data = 16'b0000100001000000;
				18'b001101111000110100: oled_data = 16'b0010000011000010;
				18'b001101111010110100: oled_data = 16'b0100000111000110;
				18'b001101111100110100: oled_data = 16'b0010000010000001;
				18'b001101111110110100: oled_data = 16'b0111000101100101;
				18'b001110000000110100: oled_data = 16'b1011101001001001;
				18'b001110000010110100: oled_data = 16'b1011001011001011;
				18'b001110000100110100: oled_data = 16'b1010101000001000;
				18'b001110000110110100: oled_data = 16'b1010101000001000;
				18'b001110001000110100: oled_data = 16'b1010101000001000;
				18'b001110001010110100: oled_data = 16'b1010101000001000;
				18'b001110001100110100: oled_data = 16'b1010101000001000;
				18'b001110001110110100: oled_data = 16'b1010101000001000;
				18'b001110010000110100: oled_data = 16'b1001000111001000;
				18'b001110010010110100: oled_data = 16'b1011010100010100;
				18'b001110010100110100: oled_data = 16'b1010111000111001;
				18'b001110010110110100: oled_data = 16'b1000110110010111;
				18'b001110011000110100: oled_data = 16'b1000110110010111;
				18'b001110011010110100: oled_data = 16'b1001110101010110;
				18'b001110011100110100: oled_data = 16'b1001101011101100;
				18'b001110011110110100: oled_data = 16'b1010000111000111;
				18'b001110100000110100: oled_data = 16'b1010000111000111;
				18'b001110100010110100: oled_data = 16'b1001100111000111;
				18'b001110100100110100: oled_data = 16'b1001100110100111;
				18'b001110100110110100: oled_data = 16'b1001100110100111;
				18'b001100011000110101: oled_data = 16'b0011000110000110;
				18'b001100011010110101: oled_data = 16'b1000101011101110;
				18'b001100011100110101: oled_data = 16'b1100101111110011;
				18'b001100011110110101: oled_data = 16'b1100001111110010;
				18'b001100100000110101: oled_data = 16'b1011101110110001;
				18'b001100100010110101: oled_data = 16'b1011101110110001;
				18'b001100100100110101: oled_data = 16'b1100001111110010;
				18'b001100100110110101: oled_data = 16'b1100001111010010;
				18'b001100101000110101: oled_data = 16'b1010001011001110;
				18'b001100101010110101: oled_data = 16'b1010001010101110;
				18'b001100101100110101: oled_data = 16'b1001001001101100;
				18'b001100101110110101: oled_data = 16'b1001101010101100;
				18'b001100110000110101: oled_data = 16'b1010101100101110;
				18'b001100110010110101: oled_data = 16'b1010101101001111;
				18'b001100110100110101: oled_data = 16'b1011001110110000;
				18'b001100110110110101: oled_data = 16'b1100010000110010;
				18'b001100111000110101: oled_data = 16'b1100110010010011;
				18'b001100111010110101: oled_data = 16'b1101010010010011;
				18'b001100111100110101: oled_data = 16'b1101010010010011;
				18'b001100111110110101: oled_data = 16'b1101010010010011;
				18'b001101000000110101: oled_data = 16'b1100010000110001;
				18'b001101000010110101: oled_data = 16'b1011001110010000;
				18'b001101000100110101: oled_data = 16'b1010101111110001;
				18'b001101000110110101: oled_data = 16'b1101111001111000;
				18'b001101001000110101: oled_data = 16'b1101111010011000;
				18'b001101001010110101: oled_data = 16'b1101111010011000;
				18'b001101001100110101: oled_data = 16'b1101111010011000;
				18'b001101001110110101: oled_data = 16'b1101111010111001;
				18'b001101010000110101: oled_data = 16'b1101011001010111;
				18'b001101010010110101: oled_data = 16'b1011110000110001;
				18'b001101010100110101: oled_data = 16'b1011110000010001;
				18'b001101010110110101: oled_data = 16'b1100110001010010;
				18'b001101011000110101: oled_data = 16'b1101010010010011;
				18'b001101011010110101: oled_data = 16'b1101010010110011;
				18'b001101011100110101: oled_data = 16'b1101010010110011;
				18'b001101011110110101: oled_data = 16'b1101010010110011;
				18'b001101100000110101: oled_data = 16'b1100010001110010;
				18'b001101100010110101: oled_data = 16'b1100110010010011;
				18'b001101100100110101: oled_data = 16'b1101010010110011;
				18'b001101100110110101: oled_data = 16'b1101010010110011;
				18'b001101101000110101: oled_data = 16'b1101010010110011;
				18'b001101101010110101: oled_data = 16'b1101010010110100;
				18'b001101101100110101: oled_data = 16'b1101010010110100;
				18'b001101101110110101: oled_data = 16'b1101010010010100;
				18'b001101110000110101: oled_data = 16'b1101010010110100;
				18'b001101110010110101: oled_data = 16'b1001001100101101;
				18'b001101110100110101: oled_data = 16'b0001000010000001;
				18'b001101110110110101: oled_data = 16'b0001000010000001;
				18'b001101111000110101: oled_data = 16'b0001100010000010;
				18'b001101111010110101: oled_data = 16'b0010000010000010;
				18'b001101111100110101: oled_data = 16'b0100000101000011;
				18'b001101111110110101: oled_data = 16'b1000000111000110;
				18'b001110000000110101: oled_data = 16'b1011001000001001;
				18'b001110000010110101: oled_data = 16'b1011001010001010;
				18'b001110000100110101: oled_data = 16'b1010100111101000;
				18'b001110000110110101: oled_data = 16'b1010101000001000;
				18'b001110001000110101: oled_data = 16'b1010101000001000;
				18'b001110001010110101: oled_data = 16'b1010101000001000;
				18'b001110001100110101: oled_data = 16'b1010100111101000;
				18'b001110001110110101: oled_data = 16'b1010000111101000;
				18'b001110010000110101: oled_data = 16'b1000100101100101;
				18'b001110010010110101: oled_data = 16'b1010001000001000;
				18'b001110010100110101: oled_data = 16'b1011001101101110;
				18'b001110010110110101: oled_data = 16'b1010010000010000;
				18'b001110011000110101: oled_data = 16'b1010001101101110;
				18'b001110011010110101: oled_data = 16'b1010001001001010;
				18'b001110011100110101: oled_data = 16'b1010000111000111;
				18'b001110011110110101: oled_data = 16'b1010000110100111;
				18'b001110100000110101: oled_data = 16'b1001100110100111;
				18'b001110100010110101: oled_data = 16'b1001100110100111;
				18'b001110100100110101: oled_data = 16'b1001100110100111;
				18'b001110100110110101: oled_data = 16'b1001100110100111;
				18'b001100011000110110: oled_data = 16'b0010100110000110;
				18'b001100011010110110: oled_data = 16'b0111001001001011;
				18'b001100011100110110: oled_data = 16'b1100001111010010;
				18'b001100011110110110: oled_data = 16'b1100001111010010;
				18'b001100100000110110: oled_data = 16'b1100001111010010;
				18'b001100100010110110: oled_data = 16'b1011001101010000;
				18'b001100100100110110: oled_data = 16'b1011101110110001;
				18'b001100100110110110: oled_data = 16'b1100001111110010;
				18'b001100101000110110: oled_data = 16'b1100001111010010;
				18'b001100101010110110: oled_data = 16'b1010101100110000;
				18'b001100101100110110: oled_data = 16'b1000101000001011;
				18'b001100101110110110: oled_data = 16'b1001001010001100;
				18'b001100110000110110: oled_data = 16'b1011001101001111;
				18'b001100110010110110: oled_data = 16'b1100010000010010;
				18'b001100110100110110: oled_data = 16'b1100110001010011;
				18'b001100110110110110: oled_data = 16'b1100110001010011;
				18'b001100111000110110: oled_data = 16'b1100110001010011;
				18'b001100111010110110: oled_data = 16'b1100110001110011;
				18'b001100111100110110: oled_data = 16'b1100110001010011;
				18'b001100111110110110: oled_data = 16'b1100010000110010;
				18'b001101000000110110: oled_data = 16'b1100010000110001;
				18'b001101000010110110: oled_data = 16'b1011110001010010;
				18'b001101000100110110: oled_data = 16'b1100110111110111;
				18'b001101000110110110: oled_data = 16'b1101011010011000;
				18'b001101001000110110: oled_data = 16'b1101011001111000;
				18'b001101001010110110: oled_data = 16'b1101011001111000;
				18'b001101001100110110: oled_data = 16'b1101011001111000;
				18'b001101001110110110: oled_data = 16'b1101011001111000;
				18'b001101010000110110: oled_data = 16'b1101111010011000;
				18'b001101010010110110: oled_data = 16'b1100010101010100;
				18'b001101010100110110: oled_data = 16'b1100010001110010;
				18'b001101010110110110: oled_data = 16'b1100110001110011;
				18'b001101011000110110: oled_data = 16'b1100110010010011;
				18'b001101011010110110: oled_data = 16'b1100110010010011;
				18'b001101011100110110: oled_data = 16'b1100110010010011;
				18'b001101011110110110: oled_data = 16'b1100110010010011;
				18'b001101100000110110: oled_data = 16'b1100010001010010;
				18'b001101100010110110: oled_data = 16'b1100110001110010;
				18'b001101100100110110: oled_data = 16'b1100110010010011;
				18'b001101100110110110: oled_data = 16'b1100110010010011;
				18'b001101101000110110: oled_data = 16'b1100110010010011;
				18'b001101101010110110: oled_data = 16'b1100110010010011;
				18'b001101101100110110: oled_data = 16'b1100110010010011;
				18'b001101101110110110: oled_data = 16'b1100110001110011;
				18'b001101110000110110: oled_data = 16'b1100110010010011;
				18'b001101110010110110: oled_data = 16'b0101100110100111;
				18'b001101110100110110: oled_data = 16'b0001100010000001;
				18'b001101110110110110: oled_data = 16'b0010100011000010;
				18'b001101111000110110: oled_data = 16'b0011100100000011;
				18'b001101111010110110: oled_data = 16'b0101100111000101;
				18'b001101111100110110: oled_data = 16'b0111001010001000;
				18'b001101111110110110: oled_data = 16'b1000101000100111;
				18'b001110000000110110: oled_data = 16'b1011001000001000;
				18'b001110000010110110: oled_data = 16'b1010101001001001;
				18'b001110000100110110: oled_data = 16'b1010100111101000;
				18'b001110000110110110: oled_data = 16'b1010100111101000;
				18'b001110001000110110: oled_data = 16'b1010100111101000;
				18'b001110001010110110: oled_data = 16'b1010000111101000;
				18'b001110001100110110: oled_data = 16'b1010100111100111;
				18'b001110001110110110: oled_data = 16'b1001100111000111;
				18'b001110010000110110: oled_data = 16'b1000100110000110;
				18'b001110010010110110: oled_data = 16'b1010000111001000;
				18'b001110010100110110: oled_data = 16'b1010000110100111;
				18'b001110010110110110: oled_data = 16'b1010000110100111;
				18'b001110011000110110: oled_data = 16'b1001100110100111;
				18'b001110011010110110: oled_data = 16'b1010000111000111;
				18'b001110011100110110: oled_data = 16'b1001100111000111;
				18'b001110011110110110: oled_data = 16'b1001100110100111;
				18'b001110100000110110: oled_data = 16'b1001100110100111;
				18'b001110100010110110: oled_data = 16'b1001100110100110;
				18'b001110100100110110: oled_data = 16'b1001000110000110;
				18'b001110100110110110: oled_data = 16'b1001000110000110;
				18'b001100011000110111: oled_data = 16'b0010100101000101;
				18'b001100011010110111: oled_data = 16'b1000001010101100;
				18'b001100011100110111: oled_data = 16'b1011101110010001;
				18'b001100011110110111: oled_data = 16'b1100001110110001;
				18'b001100100000110111: oled_data = 16'b1100001110110001;
				18'b001100100010110111: oled_data = 16'b1010101100101111;
				18'b001100100100110111: oled_data = 16'b1011001101110000;
				18'b001100100110110111: oled_data = 16'b1011101110110001;
				18'b001100101000110111: oled_data = 16'b1011101110110001;
				18'b001100101010110111: oled_data = 16'b1011101110110001;
				18'b001100101100110111: oled_data = 16'b1011001101010000;
				18'b001100101110110111: oled_data = 16'b1001101010101101;
				18'b001100110000110111: oled_data = 16'b1011001110010000;
				18'b001100110010110111: oled_data = 16'b1100001111010010;
				18'b001100110100110111: oled_data = 16'b1100101111110010;
				18'b001100110110110111: oled_data = 16'b1100110000010011;
				18'b001100111000110111: oled_data = 16'b1100110000010011;
				18'b001100111010110111: oled_data = 16'b1100110000010011;
				18'b001100111100110111: oled_data = 16'b1100001111010010;
				18'b001100111110110111: oled_data = 16'b1100001111110010;
				18'b001101000000110111: oled_data = 16'b1100010000110010;
				18'b001101000010110111: oled_data = 16'b1011010011110011;
				18'b001101000100110111: oled_data = 16'b1101011001111000;
				18'b001101000110110111: oled_data = 16'b1101011001011000;
				18'b001101001000110111: oled_data = 16'b1101011001010111;
				18'b001101001010110111: oled_data = 16'b1101011001011000;
				18'b001101001100110111: oled_data = 16'b1100111000010110;
				18'b001101001110110111: oled_data = 16'b1100010110110101;
				18'b001101010000110111: oled_data = 16'b1100111000110111;
				18'b001101010010110111: oled_data = 16'b1100010110010101;
				18'b001101010100110111: oled_data = 16'b1100010001110010;
				18'b001101010110110111: oled_data = 16'b1100110001110010;
				18'b001101011000110111: oled_data = 16'b1100110001110010;
				18'b001101011010110111: oled_data = 16'b1100110001110010;
				18'b001101011100110111: oled_data = 16'b1100110001110010;
				18'b001101011110110111: oled_data = 16'b1100110001110010;
				18'b001101100000110111: oled_data = 16'b1100010000110001;
				18'b001101100010110111: oled_data = 16'b1100110001010010;
				18'b001101100100110111: oled_data = 16'b1100110001110010;
				18'b001101100110110111: oled_data = 16'b1100110001110010;
				18'b001101101000110111: oled_data = 16'b1100110001110011;
				18'b001101101010110111: oled_data = 16'b1100110001010011;
				18'b001101101100110111: oled_data = 16'b1100110001010011;
				18'b001101101110110111: oled_data = 16'b1100110001110011;
				18'b001101110000110111: oled_data = 16'b1011001111010000;
				18'b001101110010110111: oled_data = 16'b0011000010100011;
				18'b001101110100110111: oled_data = 16'b0011100011100010;
				18'b001101110110110111: oled_data = 16'b0101000110000100;
				18'b001101111000110111: oled_data = 16'b0110101001000111;
				18'b001101111010110111: oled_data = 16'b0111101001100111;
				18'b001101111100110111: oled_data = 16'b1000001001100111;
				18'b001101111110110111: oled_data = 16'b1000101000000110;
				18'b001110000000110111: oled_data = 16'b1010100111101000;
				18'b001110000010110111: oled_data = 16'b1010001000101000;
				18'b001110000100110111: oled_data = 16'b1010100111101000;
				18'b001110000110110111: oled_data = 16'b1010100111100111;
				18'b001110001000110111: oled_data = 16'b1010000111100111;
				18'b001110001010110111: oled_data = 16'b1010000111100111;
				18'b001110001100110111: oled_data = 16'b1010000111000111;
				18'b001110001110110111: oled_data = 16'b1001100110100111;
				18'b001110010000110111: oled_data = 16'b1000100110000111;
				18'b001110010010110111: oled_data = 16'b1010000111001000;
				18'b001110010100110111: oled_data = 16'b1010000111000111;
				18'b001110010110110111: oled_data = 16'b1001100110100111;
				18'b001110011000110111: oled_data = 16'b1001000110100110;
				18'b001110011010110111: oled_data = 16'b1001100110100111;
				18'b001110011100110111: oled_data = 16'b1001100110100111;
				18'b001110011110110111: oled_data = 16'b1001100110100110;
				18'b001110100000110111: oled_data = 16'b1001100110000110;
				18'b001110100010110111: oled_data = 16'b1001000110000110;
				18'b001110100100110111: oled_data = 16'b1001000110000110;
				18'b001110100110110111: oled_data = 16'b1001000110000110;
				18'b010000011000001000: oled_data = 16'b1001101111101011;
				18'b010000011010001000: oled_data = 16'b1010010000001011;
				18'b010000011100001000: oled_data = 16'b1010010000101011;
				18'b010000011110001000: oled_data = 16'b1010110001001100;
				18'b010000100000001000: oled_data = 16'b1010110000101100;
				18'b010000100010001000: oled_data = 16'b1010110001001011;
				18'b010000100100001000: oled_data = 16'b1010110001001011;
				18'b010000100110001000: oled_data = 16'b1010110000101011;
				18'b010000101000001000: oled_data = 16'b1010110000001100;
				18'b010000101010001000: oled_data = 16'b1110011000010111;
				18'b010000101100001000: oled_data = 16'b1110110110111000;
				18'b010000101110001000: oled_data = 16'b1101110010110101;
				18'b010000110000001000: oled_data = 16'b1101110011010101;
				18'b010000110010001000: oled_data = 16'b1101110011010101;
				18'b010000110100001000: oled_data = 16'b1101110011010101;
				18'b010000110110001000: oled_data = 16'b1101110011010101;
				18'b010000111000001000: oled_data = 16'b1101110011010101;
				18'b010000111010001000: oled_data = 16'b1101110011010101;
				18'b010000111100001000: oled_data = 16'b1101110011010101;
				18'b010000111110001000: oled_data = 16'b1101110011010101;
				18'b010001000000001000: oled_data = 16'b1101110011010101;
				18'b010001000010001000: oled_data = 16'b1101110011010101;
				18'b010001000100001000: oled_data = 16'b1101110011010101;
				18'b010001000110001000: oled_data = 16'b1101110011010101;
				18'b010001001000001000: oled_data = 16'b1101110011010101;
				18'b010001001010001000: oled_data = 16'b1101110011010101;
				18'b010001001100001000: oled_data = 16'b1101110011010101;
				18'b010001001110001000: oled_data = 16'b1101110011010101;
				18'b010001010000001000: oled_data = 16'b1101110011010101;
				18'b010001010010001000: oled_data = 16'b1101110011010101;
				18'b010001010100001000: oled_data = 16'b1101110011010101;
				18'b010001010110001000: oled_data = 16'b1101110011010101;
				18'b010001011000001000: oled_data = 16'b1101110011010101;
				18'b010001011010001000: oled_data = 16'b1101110011010101;
				18'b010001011100001000: oled_data = 16'b1101110011010101;
				18'b010001011110001000: oled_data = 16'b1101110011010101;
				18'b010001100000001000: oled_data = 16'b1101110011010101;
				18'b010001100010001000: oled_data = 16'b1101110011010101;
				18'b010001100100001000: oled_data = 16'b1101110011010101;
				18'b010001100110001000: oled_data = 16'b1101110011010101;
				18'b010001101000001000: oled_data = 16'b1101010010010100;
				18'b010001101010001000: oled_data = 16'b1101110010110101;
				18'b010001101100001000: oled_data = 16'b1101110011010110;
				18'b010001101110001000: oled_data = 16'b1110010011010110;
				18'b010001110000001000: oled_data = 16'b1110010011010110;
				18'b010001110010001000: oled_data = 16'b1101110011010101;
				18'b010001110100001000: oled_data = 16'b1110010011010110;
				18'b010001110110001000: oled_data = 16'b1101110011010110;
				18'b010001111000001000: oled_data = 16'b1101110011010101;
				18'b010001111010001000: oled_data = 16'b1101110010110101;
				18'b010001111100001000: oled_data = 16'b1101010001110100;
				18'b010001111110001000: oled_data = 16'b1101110011010101;
				18'b010010000000001000: oled_data = 16'b1101110011010101;
				18'b010010000010001000: oled_data = 16'b1110010011010110;
				18'b010010000100001000: oled_data = 16'b1101110011010101;
				18'b010010000110001000: oled_data = 16'b1110111001011010;
				18'b010010001000001000: oled_data = 16'b1110011000111001;
				18'b010010001010001000: oled_data = 16'b0111001010100111;
				18'b010010001100001000: oled_data = 16'b0111001010100110;
				18'b010010001110001000: oled_data = 16'b0111101011100111;
				18'b010010010000001000: oled_data = 16'b0111101100000111;
				18'b010010010010001000: oled_data = 16'b0111101100000111;
				18'b010010010100001000: oled_data = 16'b0111001100001000;
				18'b010010010110001000: oled_data = 16'b0111001011101000;
				18'b010010011000001000: oled_data = 16'b0110101011101000;
				18'b010010011010001000: oled_data = 16'b0110001011001000;
				18'b010010011100001000: oled_data = 16'b0110001010101000;
				18'b010010011110001000: oled_data = 16'b0101101010001000;
				18'b010010100000001000: oled_data = 16'b0101101010001000;
				18'b010010100010001000: oled_data = 16'b0101001001101000;
				18'b010010100100001000: oled_data = 16'b0101001001001000;
				18'b010010100110001000: oled_data = 16'b0101001001101000;
				18'b010000011000001001: oled_data = 16'b1011010001101011;
				18'b010000011010001001: oled_data = 16'b1011010001101011;
				18'b010000011100001001: oled_data = 16'b1011010001001011;
				18'b010000011110001001: oled_data = 16'b1011010001001011;
				18'b010000100000001001: oled_data = 16'b1010110000101011;
				18'b010000100010001001: oled_data = 16'b1010110001001011;
				18'b010000100100001001: oled_data = 16'b1010110001001011;
				18'b010000100110001001: oled_data = 16'b1010110000101011;
				18'b010000101000001001: oled_data = 16'b1100010100010010;
				18'b010000101010001001: oled_data = 16'b1111011001011010;
				18'b010000101100001001: oled_data = 16'b1101110011110110;
				18'b010000101110001001: oled_data = 16'b1101110011010101;
				18'b010000110000001001: oled_data = 16'b1101010010010100;
				18'b010000110010001001: oled_data = 16'b1101110011010101;
				18'b010000110100001001: oled_data = 16'b1101110011010101;
				18'b010000110110001001: oled_data = 16'b1101110011010101;
				18'b010000111000001001: oled_data = 16'b1101110011010101;
				18'b010000111010001001: oled_data = 16'b1101110011010101;
				18'b010000111100001001: oled_data = 16'b1101110011010101;
				18'b010000111110001001: oled_data = 16'b1101110011010101;
				18'b010001000000001001: oled_data = 16'b1101110011010101;
				18'b010001000010001001: oled_data = 16'b1101110011010101;
				18'b010001000100001001: oled_data = 16'b1101110011010101;
				18'b010001000110001001: oled_data = 16'b1101110011010101;
				18'b010001001000001001: oled_data = 16'b1101110011010101;
				18'b010001001010001001: oled_data = 16'b1101110011010101;
				18'b010001001100001001: oled_data = 16'b1101110011010101;
				18'b010001001110001001: oled_data = 16'b1101110011010101;
				18'b010001010000001001: oled_data = 16'b1101110011010101;
				18'b010001010010001001: oled_data = 16'b1101110011010101;
				18'b010001010100001001: oled_data = 16'b1101110011010101;
				18'b010001010110001001: oled_data = 16'b1101110011010101;
				18'b010001011000001001: oled_data = 16'b1101110011010101;
				18'b010001011010001001: oled_data = 16'b1101110011010101;
				18'b010001011100001001: oled_data = 16'b1101110010110101;
				18'b010001011110001001: oled_data = 16'b1101010001110100;
				18'b010001100000001001: oled_data = 16'b1101110010110101;
				18'b010001100010001001: oled_data = 16'b1101110011010101;
				18'b010001100100001001: oled_data = 16'b1101110011010101;
				18'b010001100110001001: oled_data = 16'b1101110011010101;
				18'b010001101000001001: oled_data = 16'b1101110011010110;
				18'b010001101010001001: oled_data = 16'b1101110010010101;
				18'b010001101100001001: oled_data = 16'b1101010010010100;
				18'b010001101110001001: oled_data = 16'b1110010011010110;
				18'b010001110000001001: oled_data = 16'b1110010011010110;
				18'b010001110010001001: oled_data = 16'b1101110011010101;
				18'b010001110100001001: oled_data = 16'b1110010011010110;
				18'b010001110110001001: oled_data = 16'b1101110011010110;
				18'b010001111000001001: oled_data = 16'b1101110011010101;
				18'b010001111010001001: oled_data = 16'b1101110011010110;
				18'b010001111100001001: oled_data = 16'b1101010010010101;
				18'b010001111110001001: oled_data = 16'b1101110010110101;
				18'b010010000000001001: oled_data = 16'b1101110011010110;
				18'b010010000010001001: oled_data = 16'b1101110011010110;
				18'b010010000100001001: oled_data = 16'b1101110010110101;
				18'b010010000110001001: oled_data = 16'b1101110100110110;
				18'b010010001000001001: oled_data = 16'b1111011010111100;
				18'b010010001010001001: oled_data = 16'b1001101111101110;
				18'b010010001100001001: oled_data = 16'b0110101010100110;
				18'b010010001110001001: oled_data = 16'b0111101011100111;
				18'b010010010000001001: oled_data = 16'b0111101100000111;
				18'b010010010010001001: oled_data = 16'b1000001100101000;
				18'b010010010100001001: oled_data = 16'b1000001100101000;
				18'b010010010110001001: oled_data = 16'b1000101101001000;
				18'b010010011000001001: oled_data = 16'b1000101101101000;
				18'b010010011010001001: oled_data = 16'b1000101101101000;
				18'b010010011100001001: oled_data = 16'b1000101101101000;
				18'b010010011110001001: oled_data = 16'b1000101110001001;
				18'b010010100000001001: oled_data = 16'b1000101110001010;
				18'b010010100010001001: oled_data = 16'b0101101010101000;
				18'b010010100100001001: oled_data = 16'b0011101000000111;
				18'b010010100110001001: oled_data = 16'b0100001000101000;
				18'b010000011000001010: oled_data = 16'b1011010001101100;
				18'b010000011010001010: oled_data = 16'b1011010001101011;
				18'b010000011100001010: oled_data = 16'b1011010001101011;
				18'b010000011110001010: oled_data = 16'b1011010001001011;
				18'b010000100000001010: oled_data = 16'b1010110000101011;
				18'b010000100010001010: oled_data = 16'b1010010000001011;
				18'b010000100100001010: oled_data = 16'b1001001111001010;
				18'b010000100110001010: oled_data = 16'b1001001111001011;
				18'b010000101000001010: oled_data = 16'b1110011001111001;
				18'b010000101010001010: oled_data = 16'b1110010101010111;
				18'b010000101100001010: oled_data = 16'b1110010011010101;
				18'b010000101110001010: oled_data = 16'b1101010010010100;
				18'b010000110000001010: oled_data = 16'b1101110010110101;
				18'b010000110010001010: oled_data = 16'b1101110011010101;
				18'b010000110100001010: oled_data = 16'b1101110011010101;
				18'b010000110110001010: oled_data = 16'b1101110011010101;
				18'b010000111000001010: oled_data = 16'b1101110011010101;
				18'b010000111010001010: oled_data = 16'b1101110011010101;
				18'b010000111100001010: oled_data = 16'b1101110011010101;
				18'b010000111110001010: oled_data = 16'b1101110011010101;
				18'b010001000000001010: oled_data = 16'b1101110011010101;
				18'b010001000010001010: oled_data = 16'b1101110011010101;
				18'b010001000100001010: oled_data = 16'b1101110011010101;
				18'b010001000110001010: oled_data = 16'b1101110011010101;
				18'b010001001000001010: oled_data = 16'b1101110011010101;
				18'b010001001010001010: oled_data = 16'b1101110011010101;
				18'b010001001100001010: oled_data = 16'b1101110011010101;
				18'b010001001110001010: oled_data = 16'b1101110011010101;
				18'b010001010000001010: oled_data = 16'b1101110011010101;
				18'b010001010010001010: oled_data = 16'b1101110011010101;
				18'b010001010100001010: oled_data = 16'b1101110011010101;
				18'b010001010110001010: oled_data = 16'b1101110011010101;
				18'b010001011000001010: oled_data = 16'b1101110011010101;
				18'b010001011010001010: oled_data = 16'b1101110011010101;
				18'b010001011100001010: oled_data = 16'b1101110011010110;
				18'b010001011110001010: oled_data = 16'b1101110010110101;
				18'b010001100000001010: oled_data = 16'b1101010001110100;
				18'b010001100010001010: oled_data = 16'b1101110010110101;
				18'b010001100100001010: oled_data = 16'b1101110011010101;
				18'b010001100110001010: oled_data = 16'b1101110011010101;
				18'b010001101000001010: oled_data = 16'b1110010011010110;
				18'b010001101010001010: oled_data = 16'b1101110011010110;
				18'b010001101100001010: oled_data = 16'b1101010010010100;
				18'b010001101110001010: oled_data = 16'b1101010001010100;
				18'b010001110000001010: oled_data = 16'b1101110011010101;
				18'b010001110010001010: oled_data = 16'b1101110011010101;
				18'b010001110100001010: oled_data = 16'b1110010011010110;
				18'b010001110110001010: oled_data = 16'b1110010011010110;
				18'b010001111000001010: oled_data = 16'b1101110011010101;
				18'b010001111010001010: oled_data = 16'b1101110011010101;
				18'b010001111100001010: oled_data = 16'b1101110011010110;
				18'b010001111110001010: oled_data = 16'b1101010001110100;
				18'b010010000000001010: oled_data = 16'b1101110010110101;
				18'b010010000010001010: oled_data = 16'b1101110011010110;
				18'b010010000100001010: oled_data = 16'b1101110011110110;
				18'b010010000110001010: oled_data = 16'b1101010010010100;
				18'b010010001000001010: oled_data = 16'b1110010111111001;
				18'b010010001010001010: oled_data = 16'b1100110111010111;
				18'b010010001100001010: oled_data = 16'b0100100111100110;
				18'b010010001110001010: oled_data = 16'b0100101000000110;
				18'b010010010000001010: oled_data = 16'b0101101001000111;
				18'b010010010010001010: oled_data = 16'b0110101010101000;
				18'b010010010100001010: oled_data = 16'b0111101011101000;
				18'b010010010110001010: oled_data = 16'b1000001100100111;
				18'b010010011000001010: oled_data = 16'b1000101101001000;
				18'b010010011010001010: oled_data = 16'b1000101101101000;
				18'b010010011100001010: oled_data = 16'b1000101110001000;
				18'b010010011110001010: oled_data = 16'b1000101110001000;
				18'b010010100000001010: oled_data = 16'b1000101110001001;
				18'b010010100010001010: oled_data = 16'b0111001011101001;
				18'b010010100100001010: oled_data = 16'b1001001101001101;
				18'b010010100110001010: oled_data = 16'b1011010000110001;
				18'b010000011000001011: oled_data = 16'b1001001111001010;
				18'b010000011010001011: oled_data = 16'b1000101110001010;
				18'b010000011100001011: oled_data = 16'b0111101100101001;
				18'b010000011110001011: oled_data = 16'b0111001011101001;
				18'b010000100000001011: oled_data = 16'b0110001010101000;
				18'b010000100010001011: oled_data = 16'b0110001010001000;
				18'b010000100100001011: oled_data = 16'b0101101001101000;
				18'b010000100110001011: oled_data = 16'b1001110001010000;
				18'b010000101000001011: oled_data = 16'b1110111000111010;
				18'b010000101010001011: oled_data = 16'b1101110011110110;
				18'b010000101100001011: oled_data = 16'b1101110010110101;
				18'b010000101110001011: oled_data = 16'b1101110010010100;
				18'b010000110000001011: oled_data = 16'b1101110011010110;
				18'b010000110010001011: oled_data = 16'b1101110011010101;
				18'b010000110100001011: oled_data = 16'b1101110011010101;
				18'b010000110110001011: oled_data = 16'b1101110011010101;
				18'b010000111000001011: oled_data = 16'b1101110011010101;
				18'b010000111010001011: oled_data = 16'b1101110011010101;
				18'b010000111100001011: oled_data = 16'b1101110011010101;
				18'b010000111110001011: oled_data = 16'b1101110011010101;
				18'b010001000000001011: oled_data = 16'b1101110011010101;
				18'b010001000010001011: oled_data = 16'b1101110011010101;
				18'b010001000100001011: oled_data = 16'b1101110011010101;
				18'b010001000110001011: oled_data = 16'b1101110011010101;
				18'b010001001000001011: oled_data = 16'b1101110011010101;
				18'b010001001010001011: oled_data = 16'b1101110011010101;
				18'b010001001100001011: oled_data = 16'b1101110011010101;
				18'b010001001110001011: oled_data = 16'b1101110011010101;
				18'b010001010000001011: oled_data = 16'b1101110011010101;
				18'b010001010010001011: oled_data = 16'b1101110011010101;
				18'b010001010100001011: oled_data = 16'b1101110011010101;
				18'b010001010110001011: oled_data = 16'b1101110011010101;
				18'b010001011000001011: oled_data = 16'b1101110011010101;
				18'b010001011010001011: oled_data = 16'b1101110011010101;
				18'b010001011100001011: oled_data = 16'b1101110011010101;
				18'b010001011110001011: oled_data = 16'b1101110011010101;
				18'b010001100000001011: oled_data = 16'b1101110011010101;
				18'b010001100010001011: oled_data = 16'b1101010001110100;
				18'b010001100100001011: oled_data = 16'b1101110010110101;
				18'b010001100110001011: oled_data = 16'b1101110011010101;
				18'b010001101000001011: oled_data = 16'b1110010100110110;
				18'b010001101010001011: oled_data = 16'b1110010100010110;
				18'b010001101100001011: oled_data = 16'b1101110011010110;
				18'b010001101110001011: oled_data = 16'b1100110000110011;
				18'b010001110000001011: oled_data = 16'b1100001111110010;
				18'b010001110010001011: oled_data = 16'b1101110011010110;
				18'b010001110100001011: oled_data = 16'b1110010011010110;
				18'b010001110110001011: oled_data = 16'b1101110011010101;
				18'b010001111000001011: oled_data = 16'b1101110011010101;
				18'b010001111010001011: oled_data = 16'b1101110011010101;
				18'b010001111100001011: oled_data = 16'b1101110011010110;
				18'b010001111110001011: oled_data = 16'b1101110010110101;
				18'b010010000000001011: oled_data = 16'b1101010010010101;
				18'b010010000010001011: oled_data = 16'b1101110011010110;
				18'b010010000100001011: oled_data = 16'b1101110011110110;
				18'b010010000110001011: oled_data = 16'b1101110010110101;
				18'b010010001000001011: oled_data = 16'b1101110011110110;
				18'b010010001010001011: oled_data = 16'b1110111001111010;
				18'b010010001100001011: oled_data = 16'b0100101001001000;
				18'b010010001110001011: oled_data = 16'b0010000100100101;
				18'b010010010000001011: oled_data = 16'b0010100101000101;
				18'b010010010010001011: oled_data = 16'b0011000110000110;
				18'b010010010100001011: oled_data = 16'b0011100111000111;
				18'b010010010110001011: oled_data = 16'b0100001000000110;
				18'b010010011000001011: oled_data = 16'b0101001000100111;
				18'b010010011010001011: oled_data = 16'b0101101001100111;
				18'b010010011100001011: oled_data = 16'b0111001011001000;
				18'b010010011110001011: oled_data = 16'b1010001110001100;
				18'b010010100000001011: oled_data = 16'b1100010001010000;
				18'b010010100010001011: oled_data = 16'b1101110010110010;
				18'b010010100100001011: oled_data = 16'b1101110001010001;
				18'b010010100110001011: oled_data = 16'b1100101110001110;
				18'b010000011000001100: oled_data = 16'b0110001010101000;
				18'b010000011010001100: oled_data = 16'b0110001010101000;
				18'b010000011100001100: oled_data = 16'b0110101011101001;
				18'b010000011110001100: oled_data = 16'b0111101100101010;
				18'b010000100000001100: oled_data = 16'b1000001101001010;
				18'b010000100010001100: oled_data = 16'b1001001110001010;
				18'b010000100100001100: oled_data = 16'b1001101111001011;
				18'b010000100110001100: oled_data = 16'b1101110111110111;
				18'b010000101000001100: oled_data = 16'b1110010101010111;
				18'b010000101010001100: oled_data = 16'b1110010011010110;
				18'b010000101100001100: oled_data = 16'b1101110010010101;
				18'b010000101110001100: oled_data = 16'b1101110010110101;
				18'b010000110000001100: oled_data = 16'b1101110011010101;
				18'b010000110010001100: oled_data = 16'b1101110011010101;
				18'b010000110100001100: oled_data = 16'b1101110011010101;
				18'b010000110110001100: oled_data = 16'b1101110011010101;
				18'b010000111000001100: oled_data = 16'b1101110011010101;
				18'b010000111010001100: oled_data = 16'b1101110011010101;
				18'b010000111100001100: oled_data = 16'b1101110011010101;
				18'b010000111110001100: oled_data = 16'b1101110011010101;
				18'b010001000000001100: oled_data = 16'b1101110011010101;
				18'b010001000010001100: oled_data = 16'b1101110011010101;
				18'b010001000100001100: oled_data = 16'b1101110011010101;
				18'b010001000110001100: oled_data = 16'b1101110011010101;
				18'b010001001000001100: oled_data = 16'b1101110011010101;
				18'b010001001010001100: oled_data = 16'b1101110010010101;
				18'b010001001100001100: oled_data = 16'b1101110010110101;
				18'b010001001110001100: oled_data = 16'b1101110011010101;
				18'b010001010000001100: oled_data = 16'b1101110011010101;
				18'b010001010010001100: oled_data = 16'b1101110011010101;
				18'b010001010100001100: oled_data = 16'b1101110011010101;
				18'b010001010110001100: oled_data = 16'b1101110011010101;
				18'b010001011000001100: oled_data = 16'b1101110011010101;
				18'b010001011010001100: oled_data = 16'b1101110011010101;
				18'b010001011100001100: oled_data = 16'b1101110011010101;
				18'b010001011110001100: oled_data = 16'b1101110011010101;
				18'b010001100000001100: oled_data = 16'b1101110011010110;
				18'b010001100010001100: oled_data = 16'b1101110011010101;
				18'b010001100100001100: oled_data = 16'b1100110000110011;
				18'b010001100110001100: oled_data = 16'b1101110010110101;
				18'b010001101000001100: oled_data = 16'b1110010011110110;
				18'b010001101010001100: oled_data = 16'b1110110101010111;
				18'b010001101100001100: oled_data = 16'b1101110011010110;
				18'b010001101110001100: oled_data = 16'b1110010011010110;
				18'b010001110000001100: oled_data = 16'b1100001111110010;
				18'b010001110010001100: oled_data = 16'b1100001111110010;
				18'b010001110100001100: oled_data = 16'b1110010011110110;
				18'b010001110110001100: oled_data = 16'b1101110011010101;
				18'b010001111000001100: oled_data = 16'b1101110011010110;
				18'b010001111010001100: oled_data = 16'b1101110011010110;
				18'b010001111100001100: oled_data = 16'b1101110011010110;
				18'b010001111110001100: oled_data = 16'b1110010011110110;
				18'b010010000000001100: oled_data = 16'b1101010001110100;
				18'b010010000010001100: oled_data = 16'b1101110010110101;
				18'b010010000100001100: oled_data = 16'b1101110011010110;
				18'b010010000110001100: oled_data = 16'b1101110010110101;
				18'b010010001000001100: oled_data = 16'b1101010010010100;
				18'b010010001010001100: oled_data = 16'b1110110111111001;
				18'b010010001100001100: oled_data = 16'b1000101111010000;
				18'b010010001110001100: oled_data = 16'b0001100100000100;
				18'b010010010000001100: oled_data = 16'b0010000101000110;
				18'b010010010010001100: oled_data = 16'b0010100101100110;
				18'b010010010100001100: oled_data = 16'b0010100110000111;
				18'b010010010110001100: oled_data = 16'b0010100110000111;
				18'b010010011000001100: oled_data = 16'b0010100110100111;
				18'b010010011010001100: oled_data = 16'b0110101010101010;
				18'b010010011100001100: oled_data = 16'b1011110001010001;
				18'b010010011110001100: oled_data = 16'b1110010011010100;
				18'b010010100000001100: oled_data = 16'b1101110000110001;
				18'b010010100010001100: oled_data = 16'b1100001100001100;
				18'b010010100100001100: oled_data = 16'b1010101001001001;
				18'b010010100110001100: oled_data = 16'b1010101000001000;
				18'b010000011000001101: oled_data = 16'b1010010000001011;
				18'b010000011010001101: oled_data = 16'b1010010000101011;
				18'b010000011100001101: oled_data = 16'b1010010001001100;
				18'b010000011110001101: oled_data = 16'b1010110000101100;
				18'b010000100000001101: oled_data = 16'b1010110000001011;
				18'b010000100010001101: oled_data = 16'b1010110000001011;
				18'b010000100100001101: oled_data = 16'b1011010001101101;
				18'b010000100110001101: oled_data = 16'b1110110111111000;
				18'b010000101000001101: oled_data = 16'b1101110011010110;
				18'b010000101010001101: oled_data = 16'b1101110011010101;
				18'b010000101100001101: oled_data = 16'b1101010010010100;
				18'b010000101110001101: oled_data = 16'b1101110011010110;
				18'b010000110000001101: oled_data = 16'b1101110011010101;
				18'b010000110010001101: oled_data = 16'b1101110011010101;
				18'b010000110100001101: oled_data = 16'b1101110011010110;
				18'b010000110110001101: oled_data = 16'b1101110010010101;
				18'b010000111000001101: oled_data = 16'b1101110010110101;
				18'b010000111010001101: oled_data = 16'b1101110011010101;
				18'b010000111100001101: oled_data = 16'b1101110011010101;
				18'b010000111110001101: oled_data = 16'b1101110011010101;
				18'b010001000000001101: oled_data = 16'b1101110011010101;
				18'b010001000010001101: oled_data = 16'b1101110011010101;
				18'b010001000100001101: oled_data = 16'b1101110011010101;
				18'b010001000110001101: oled_data = 16'b1101110011010101;
				18'b010001001000001101: oled_data = 16'b1101110011010110;
				18'b010001001010001101: oled_data = 16'b1101010001110100;
				18'b010001001100001101: oled_data = 16'b1101110010110101;
				18'b010001001110001101: oled_data = 16'b1101110011010110;
				18'b010001010000001101: oled_data = 16'b1101110011010101;
				18'b010001010010001101: oled_data = 16'b1101110011010101;
				18'b010001010100001101: oled_data = 16'b1101110011010101;
				18'b010001010110001101: oled_data = 16'b1101110011010101;
				18'b010001011000001101: oled_data = 16'b1101110011010101;
				18'b010001011010001101: oled_data = 16'b1101110011010101;
				18'b010001011100001101: oled_data = 16'b1101110011010101;
				18'b010001011110001101: oled_data = 16'b1101110011010101;
				18'b010001100000001101: oled_data = 16'b1101110011010101;
				18'b010001100010001101: oled_data = 16'b1101110011010110;
				18'b010001100100001101: oled_data = 16'b1101010010110101;
				18'b010001100110001101: oled_data = 16'b1100110000110011;
				18'b010001101000001101: oled_data = 16'b1101110011010101;
				18'b010001101010001101: oled_data = 16'b1110010011110110;
				18'b010001101100001101: oled_data = 16'b1101110011010101;
				18'b010001101110001101: oled_data = 16'b1101110011010101;
				18'b010001110000001101: oled_data = 16'b1101110011010101;
				18'b010001110010001101: oled_data = 16'b1011101110110001;
				18'b010001110100001101: oled_data = 16'b1100110000110011;
				18'b010001110110001101: oled_data = 16'b1110010011010110;
				18'b010001111000001101: oled_data = 16'b1101110011010110;
				18'b010001111010001101: oled_data = 16'b1101110011010110;
				18'b010001111100001101: oled_data = 16'b1101110011010110;
				18'b010001111110001101: oled_data = 16'b1110010011110110;
				18'b010010000000001101: oled_data = 16'b1101110010110101;
				18'b010010000010001101: oled_data = 16'b1101010010010100;
				18'b010010000100001101: oled_data = 16'b1101110011010110;
				18'b010010000110001101: oled_data = 16'b1101110011010101;
				18'b010010001000001101: oled_data = 16'b1101010001010100;
				18'b010010001010001101: oled_data = 16'b1101110101010111;
				18'b010010001100001101: oled_data = 16'b1011010011110100;
				18'b010010001110001101: oled_data = 16'b0010000100000100;
				18'b010010010000001101: oled_data = 16'b0010000101000110;
				18'b010010010010001101: oled_data = 16'b0010000101000110;
				18'b010010010100001101: oled_data = 16'b0010000101000110;
				18'b010010010110001101: oled_data = 16'b0100001000001000;
				18'b010010011000001101: oled_data = 16'b1010101111110000;
				18'b010010011010001101: oled_data = 16'b1110010100010100;
				18'b010010011100001101: oled_data = 16'b1110010010010010;
				18'b010010011110001101: oled_data = 16'b1100001100101101;
				18'b010010100000001101: oled_data = 16'b1011001001001001;
				18'b010010100010001101: oled_data = 16'b1011001000101000;
				18'b010010100100001101: oled_data = 16'b1010101000101000;
				18'b010010100110001101: oled_data = 16'b1010101000001000;
				18'b010000011000001110: oled_data = 16'b1011010001101011;
				18'b010000011010001110: oled_data = 16'b1011010001101100;
				18'b010000011100001110: oled_data = 16'b1011010001101011;
				18'b010000011110001110: oled_data = 16'b1010110001001010;
				18'b010000100000001110: oled_data = 16'b1010110000101011;
				18'b010000100010001110: oled_data = 16'b1010010000001010;
				18'b010000100100001110: oled_data = 16'b1100010100010001;
				18'b010000100110001110: oled_data = 16'b1110010101110111;
				18'b010000101000001110: oled_data = 16'b1101110011010110;
				18'b010000101010001110: oled_data = 16'b1101010010010100;
				18'b010000101100001110: oled_data = 16'b1101110010010101;
				18'b010000101110001110: oled_data = 16'b1101110011010110;
				18'b010000110000001110: oled_data = 16'b1101110011010101;
				18'b010000110010001110: oled_data = 16'b1101110011010101;
				18'b010000110100001110: oled_data = 16'b1101110011010101;
				18'b010000110110001110: oled_data = 16'b1101010001110100;
				18'b010000111000001110: oled_data = 16'b1101110011010101;
				18'b010000111010001110: oled_data = 16'b1101110011010110;
				18'b010000111100001110: oled_data = 16'b1101110011010101;
				18'b010000111110001110: oled_data = 16'b1101110011010101;
				18'b010001000000001110: oled_data = 16'b1101110011010101;
				18'b010001000010001110: oled_data = 16'b1101110010110101;
				18'b010001000100001110: oled_data = 16'b1101010010010101;
				18'b010001000110001110: oled_data = 16'b1101110011010110;
				18'b010001001000001110: oled_data = 16'b1101110011010110;
				18'b010001001010001110: oled_data = 16'b1101110010010101;
				18'b010001001100001110: oled_data = 16'b1101010010010100;
				18'b010001001110001110: oled_data = 16'b1101110011010110;
				18'b010001010000001110: oled_data = 16'b1101110011010101;
				18'b010001010010001110: oled_data = 16'b1101110011010101;
				18'b010001010100001110: oled_data = 16'b1101110011010101;
				18'b010001010110001110: oled_data = 16'b1101110011010101;
				18'b010001011000001110: oled_data = 16'b1101110011010101;
				18'b010001011010001110: oled_data = 16'b1101110011010101;
				18'b010001011100001110: oled_data = 16'b1101110011010101;
				18'b010001011110001110: oled_data = 16'b1101110011010101;
				18'b010001100000001110: oled_data = 16'b1101110011010101;
				18'b010001100010001110: oled_data = 16'b1101110011010101;
				18'b010001100100001110: oled_data = 16'b1110010011110110;
				18'b010001100110001110: oled_data = 16'b1101010001110100;
				18'b010001101000001110: oled_data = 16'b1100110001010011;
				18'b010001101010001110: oled_data = 16'b1101010011010101;
				18'b010001101100001110: oled_data = 16'b1101110011010110;
				18'b010001101110001110: oled_data = 16'b1101110011010101;
				18'b010001110000001110: oled_data = 16'b1101110011010110;
				18'b010001110010001110: oled_data = 16'b1101010010010101;
				18'b010001110100001110: oled_data = 16'b1011001101010000;
				18'b010001110110001110: oled_data = 16'b1100110000110011;
				18'b010001111000001110: oled_data = 16'b1101110011010110;
				18'b010001111010001110: oled_data = 16'b1101110011010110;
				18'b010001111100001110: oled_data = 16'b1101110011010110;
				18'b010001111110001110: oled_data = 16'b1101110011010110;
				18'b010010000000001110: oled_data = 16'b1101110011010110;
				18'b010010000010001110: oled_data = 16'b1101010001110100;
				18'b010010000100001110: oled_data = 16'b1101110011010101;
				18'b010010000110001110: oled_data = 16'b1101110011010101;
				18'b010010001000001110: oled_data = 16'b1101010001110100;
				18'b010010001010001110: oled_data = 16'b1101110011010101;
				18'b010010001100001110: oled_data = 16'b1100010011110101;
				18'b010010001110001110: oled_data = 16'b0010100101100110;
				18'b010010010000001110: oled_data = 16'b0010000100100101;
				18'b010010010010001110: oled_data = 16'b0010000100100101;
				18'b010010010100001110: oled_data = 16'b0110001010001001;
				18'b010010010110001110: oled_data = 16'b1101010010010010;
				18'b010010011000001110: oled_data = 16'b1110110011110100;
				18'b010010011010001110: oled_data = 16'b1101001111001111;
				18'b010010011100001110: oled_data = 16'b1011001010001010;
				18'b010010011110001110: oled_data = 16'b1011001000001000;
				18'b010010100000001110: oled_data = 16'b1011001000101001;
				18'b010010100010001110: oled_data = 16'b1011001000101000;
				18'b010010100100001110: oled_data = 16'b1010101000101000;
				18'b010010100110001110: oled_data = 16'b1010101000001000;
				18'b010000011000001111: oled_data = 16'b1011010001001011;
				18'b010000011010001111: oled_data = 16'b1010110000101011;
				18'b010000011100001111: oled_data = 16'b1010010000001011;
				18'b010000011110001111: oled_data = 16'b1001001111001001;
				18'b010000100000001111: oled_data = 16'b1000001101001001;
				18'b010000100010001111: oled_data = 16'b0111101011101000;
				18'b010000100100001111: oled_data = 16'b1100110100110101;
				18'b010000100110001111: oled_data = 16'b1101110100110111;
				18'b010000101000001111: oled_data = 16'b1101110011010110;
				18'b010000101010001111: oled_data = 16'b1101010001110100;
				18'b010000101100001111: oled_data = 16'b1101110011010110;
				18'b010000101110001111: oled_data = 16'b1101110011010101;
				18'b010000110000001111: oled_data = 16'b1101110011010101;
				18'b010000110010001111: oled_data = 16'b1101110011010101;
				18'b010000110100001111: oled_data = 16'b1101110011010101;
				18'b010000110110001111: oled_data = 16'b1101010001110100;
				18'b010000111000001111: oled_data = 16'b1110010011010110;
				18'b010000111010001111: oled_data = 16'b1101110011010101;
				18'b010000111100001111: oled_data = 16'b1101110011010101;
				18'b010000111110001111: oled_data = 16'b1101110011010101;
				18'b010001000000001111: oled_data = 16'b1101110011010101;
				18'b010001000010001111: oled_data = 16'b1101110010110101;
				18'b010001000100001111: oled_data = 16'b1101010010010100;
				18'b010001000110001111: oled_data = 16'b1101110011010110;
				18'b010001001000001111: oled_data = 16'b1101110011010101;
				18'b010001001010001111: oled_data = 16'b1101110010110101;
				18'b010001001100001111: oled_data = 16'b1101010010010100;
				18'b010001001110001111: oled_data = 16'b1101110011010101;
				18'b010001010000001111: oled_data = 16'b1101110011010101;
				18'b010001010010001111: oled_data = 16'b1101110011010101;
				18'b010001010100001111: oled_data = 16'b1101110011010101;
				18'b010001010110001111: oled_data = 16'b1101110011010101;
				18'b010001011000001111: oled_data = 16'b1101110011010101;
				18'b010001011010001111: oled_data = 16'b1101110011010110;
				18'b010001011100001111: oled_data = 16'b1101110011010101;
				18'b010001011110001111: oled_data = 16'b1101110011010101;
				18'b010001100000001111: oled_data = 16'b1101110011010101;
				18'b010001100010001111: oled_data = 16'b1101110011010101;
				18'b010001100100001111: oled_data = 16'b1101110011010101;
				18'b010001100110001111: oled_data = 16'b1101110010110101;
				18'b010001101000001111: oled_data = 16'b1101010011010101;
				18'b010001101010001111: oled_data = 16'b1100110011010101;
				18'b010001101100001111: oled_data = 16'b1101010010110101;
				18'b010001101110001111: oled_data = 16'b1101110011010110;
				18'b010001110000001111: oled_data = 16'b1101110011010101;
				18'b010001110010001111: oled_data = 16'b1110010011110110;
				18'b010001110100001111: oled_data = 16'b1100001111110010;
				18'b010001110110001111: oled_data = 16'b1010101100101111;
				18'b010001111000001111: oled_data = 16'b1100110000110011;
				18'b010001111010001111: oled_data = 16'b1101110011110110;
				18'b010001111100001111: oled_data = 16'b1101110011010110;
				18'b010001111110001111: oled_data = 16'b1101110011010101;
				18'b010010000000001111: oled_data = 16'b1101110011010110;
				18'b010010000010001111: oled_data = 16'b1101010010010100;
				18'b010010000100001111: oled_data = 16'b1101110010110101;
				18'b010010000110001111: oled_data = 16'b1110010011010110;
				18'b010010001000001111: oled_data = 16'b1101010010010100;
				18'b010010001010001111: oled_data = 16'b1101110011010101;
				18'b010010001100001111: oled_data = 16'b1101010011110101;
				18'b010010001110001111: oled_data = 16'b0011100110100111;
				18'b010010010000001111: oled_data = 16'b0001100100000101;
				18'b010010010010001111: oled_data = 16'b0111101100001100;
				18'b010010010100001111: oled_data = 16'b1110010100010100;
				18'b010010010110001111: oled_data = 16'b1110010010110010;
				18'b010010011000001111: oled_data = 16'b1100001100001100;
				18'b010010011010001111: oled_data = 16'b1011001000101001;
				18'b010010011100001111: oled_data = 16'b1011001000101001;
				18'b010010011110001111: oled_data = 16'b1011001000101001;
				18'b010010100000001111: oled_data = 16'b1011001000101001;
				18'b010010100010001111: oled_data = 16'b1011001000101000;
				18'b010010100100001111: oled_data = 16'b1010101000101000;
				18'b010010100110001111: oled_data = 16'b1010101000001000;
				18'b010000011000010000: oled_data = 16'b0110101011001010;
				18'b010000011010010000: oled_data = 16'b0101101010101001;
				18'b010000011100010000: oled_data = 16'b0101001010001010;
				18'b010000011110010000: oled_data = 16'b0100001001001001;
				18'b010000100000010000: oled_data = 16'b0011101000101000;
				18'b010000100010010000: oled_data = 16'b0100001001001001;
				18'b010000100100010000: oled_data = 16'b1100110100110110;
				18'b010000100110010000: oled_data = 16'b1101110011110110;
				18'b010000101000010000: oled_data = 16'b1101110010110101;
				18'b010000101010010000: oled_data = 16'b1101010010010100;
				18'b010000101100010000: oled_data = 16'b1101110011010110;
				18'b010000101110010000: oled_data = 16'b1101110011010110;
				18'b010000110000010000: oled_data = 16'b1101110011010101;
				18'b010000110010010000: oled_data = 16'b1101110011010101;
				18'b010000110100010000: oled_data = 16'b1101110010110101;
				18'b010000110110010000: oled_data = 16'b1101110010110101;
				18'b010000111000010000: oled_data = 16'b1110010011010110;
				18'b010000111010010000: oled_data = 16'b1101110010110101;
				18'b010000111100010000: oled_data = 16'b1101110010110101;
				18'b010000111110010000: oled_data = 16'b1101110011010101;
				18'b010001000000010000: oled_data = 16'b1101110011010101;
				18'b010001000010010000: oled_data = 16'b1101110010110101;
				18'b010001000100010000: oled_data = 16'b1101010001110100;
				18'b010001000110010000: oled_data = 16'b1101110011010110;
				18'b010001001000010000: oled_data = 16'b1101110011010101;
				18'b010001001010010000: oled_data = 16'b1101110011010110;
				18'b010001001100010000: oled_data = 16'b1101110010010101;
				18'b010001001110010000: oled_data = 16'b1101110011010101;
				18'b010001010000010000: oled_data = 16'b1101110011010101;
				18'b010001010010010000: oled_data = 16'b1101110011010101;
				18'b010001010100010000: oled_data = 16'b1101110011010101;
				18'b010001010110010000: oled_data = 16'b1101110011010101;
				18'b010001011000010000: oled_data = 16'b1101110011010101;
				18'b010001011010010000: oled_data = 16'b1110110101010111;
				18'b010001011100010000: oled_data = 16'b1101110011110110;
				18'b010001011110010000: oled_data = 16'b1101110011010101;
				18'b010001100000010000: oled_data = 16'b1101110011010101;
				18'b010001100010010000: oled_data = 16'b1101110011010101;
				18'b010001100100010000: oled_data = 16'b1101110010110101;
				18'b010001100110010000: oled_data = 16'b1101110011010101;
				18'b010001101000010000: oled_data = 16'b1101110011010101;
				18'b010001101010010000: oled_data = 16'b1110010110111000;
				18'b010001101100010000: oled_data = 16'b1100110011110101;
				18'b010001101110010000: oled_data = 16'b1101110010110101;
				18'b010001110000010000: oled_data = 16'b1101110011010110;
				18'b010001110010010000: oled_data = 16'b1101110011010110;
				18'b010001110100010000: oled_data = 16'b1101110010110101;
				18'b010001110110010000: oled_data = 16'b1011101110010001;
				18'b010001111000010000: oled_data = 16'b1011001101010000;
				18'b010001111010010000: oled_data = 16'b1100110000110011;
				18'b010001111100010000: oled_data = 16'b1110010011010110;
				18'b010001111110010000: oled_data = 16'b1101110011010101;
				18'b010010000000010000: oled_data = 16'b1101110011010110;
				18'b010010000010010000: oled_data = 16'b1101110010110101;
				18'b010010000100010000: oled_data = 16'b1101110010010101;
				18'b010010000110010000: oled_data = 16'b1110010011110110;
				18'b010010001000010000: oled_data = 16'b1101010010010100;
				18'b010010001010010000: oled_data = 16'b1101110010110101;
				18'b010010001100010000: oled_data = 16'b1101010011010101;
				18'b010010001110010000: oled_data = 16'b0101101001101010;
				18'b010010010000010000: oled_data = 16'b1000001100001101;
				18'b010010010010010000: oled_data = 16'b1110110100110101;
				18'b010010010100010000: oled_data = 16'b1101110001010001;
				18'b010010010110010000: oled_data = 16'b1011101010101010;
				18'b010010011000010000: oled_data = 16'b1011001000101001;
				18'b010010011010010000: oled_data = 16'b1011001000101001;
				18'b010010011100010000: oled_data = 16'b1011001001001001;
				18'b010010011110010000: oled_data = 16'b1011001000101001;
				18'b010010100000010000: oled_data = 16'b1011001000101001;
				18'b010010100010010000: oled_data = 16'b1011001000101000;
				18'b010010100100010000: oled_data = 16'b1010101000101000;
				18'b010010100110010000: oled_data = 16'b1010101000001000;
				18'b010000011000010001: oled_data = 16'b0011101001001010;
				18'b010000011010010001: oled_data = 16'b0110010001010011;
				18'b010000011100010001: oled_data = 16'b0110010011110101;
				18'b010000011110010001: oled_data = 16'b0110010010110100;
				18'b010000100000010001: oled_data = 16'b0100101110110000;
				18'b010000100010010001: oled_data = 16'b0100101100001101;
				18'b010000100100010001: oled_data = 16'b1101010100110111;
				18'b010000100110010001: oled_data = 16'b1110010011010110;
				18'b010000101000010001: oled_data = 16'b1101110010110101;
				18'b010000101010010001: oled_data = 16'b1101010010010101;
				18'b010000101100010001: oled_data = 16'b1101110011010110;
				18'b010000101110010001: oled_data = 16'b1101110011010110;
				18'b010000110000010001: oled_data = 16'b1101110011010101;
				18'b010000110010010001: oled_data = 16'b1101110011010110;
				18'b010000110100010001: oled_data = 16'b1101110010010101;
				18'b010000110110010001: oled_data = 16'b1101110010010101;
				18'b010000111000010001: oled_data = 16'b1110010011010110;
				18'b010000111010010001: oled_data = 16'b1101010010010100;
				18'b010000111100010001: oled_data = 16'b1101110010110101;
				18'b010000111110010001: oled_data = 16'b1101110011010101;
				18'b010001000000010001: oled_data = 16'b1101110011010101;
				18'b010001000010010001: oled_data = 16'b1101110010110101;
				18'b010001000100010001: oled_data = 16'b1101010001110100;
				18'b010001000110010001: oled_data = 16'b1101110011010110;
				18'b010001001000010001: oled_data = 16'b1101110011010101;
				18'b010001001010010001: oled_data = 16'b1110010011010110;
				18'b010001001100010001: oled_data = 16'b1101010010010100;
				18'b010001001110010001: oled_data = 16'b1101110010110101;
				18'b010001010000010001: oled_data = 16'b1101110011010101;
				18'b010001010010010001: oled_data = 16'b1101110011010101;
				18'b010001010100010001: oled_data = 16'b1101110011010101;
				18'b010001010110010001: oled_data = 16'b1101110011010101;
				18'b010001011000010001: oled_data = 16'b1101110010110101;
				18'b010001011010010001: oled_data = 16'b1110010101010111;
				18'b010001011100010001: oled_data = 16'b1110110100110111;
				18'b010001011110010001: oled_data = 16'b1101110011010101;
				18'b010001100000010001: oled_data = 16'b1101110011010101;
				18'b010001100010010001: oled_data = 16'b1101110011010101;
				18'b010001100100010001: oled_data = 16'b1101110010110101;
				18'b010001100110010001: oled_data = 16'b1101010010010101;
				18'b010001101000010001: oled_data = 16'b1101110010110101;
				18'b010001101010010001: oled_data = 16'b1101010100110110;
				18'b010001101100010001: oled_data = 16'b1110011001011000;
				18'b010001101110010001: oled_data = 16'b1101010100010101;
				18'b010001110000010001: oled_data = 16'b1101110011010110;
				18'b010001110010010001: oled_data = 16'b1101110011010101;
				18'b010001110100010001: oled_data = 16'b1110010011010110;
				18'b010001110110010001: oled_data = 16'b1100001111110010;
				18'b010001111000010001: oled_data = 16'b1011001101110000;
				18'b010001111010010001: oled_data = 16'b1011001101110001;
				18'b010001111100010001: oled_data = 16'b1101010001110100;
				18'b010001111110010001: oled_data = 16'b1110010011010110;
				18'b010010000000010001: oled_data = 16'b1101110011010101;
				18'b010010000010010001: oled_data = 16'b1101110011010101;
				18'b010010000100010001: oled_data = 16'b1101010010010100;
				18'b010010000110010001: oled_data = 16'b1110010011110110;
				18'b010010001000010001: oled_data = 16'b1101010010010100;
				18'b010010001010010001: oled_data = 16'b1101110010010101;
				18'b010010001100010001: oled_data = 16'b1101010010010101;
				18'b010010001110010001: oled_data = 16'b1011110000110010;
				18'b010010010000010001: oled_data = 16'b1110010100010100;
				18'b010010010010010001: oled_data = 16'b1101010000010000;
				18'b010010010100010001: oled_data = 16'b1011001001101010;
				18'b010010010110010001: oled_data = 16'b1011001000101001;
				18'b010010011000010001: oled_data = 16'b1011001001001001;
				18'b010010011010010001: oled_data = 16'b1011001000101001;
				18'b010010011100010001: oled_data = 16'b1011001001001001;
				18'b010010011110010001: oled_data = 16'b1011001000101001;
				18'b010010100000010001: oled_data = 16'b1011001000101001;
				18'b010010100010010001: oled_data = 16'b1011001000101000;
				18'b010010100100010001: oled_data = 16'b1011001000001000;
				18'b010010100110010001: oled_data = 16'b1011001000001000;
				18'b010000011000010010: oled_data = 16'b0101001101101111;
				18'b010000011010010010: oled_data = 16'b0111111000111010;
				18'b010000011100010010: oled_data = 16'b0111111001011010;
				18'b010000011110010010: oled_data = 16'b0111111001011010;
				18'b010000100000010010: oled_data = 16'b0111111000111010;
				18'b010000100010010010: oled_data = 16'b0111111000111000;
				18'b010000100100010010: oled_data = 16'b1001110111111001;
				18'b010000100110010010: oled_data = 16'b1011110101010111;
				18'b010000101000010010: oled_data = 16'b1101010010110101;
				18'b010000101010010010: oled_data = 16'b1101110010110101;
				18'b010000101100010010: oled_data = 16'b1101110011010110;
				18'b010000101110010010: oled_data = 16'b1101110011010110;
				18'b010000110000010010: oled_data = 16'b1101110011010101;
				18'b010000110010010010: oled_data = 16'b1101110011010110;
				18'b010000110100010010: oled_data = 16'b1101010010010101;
				18'b010000110110010010: oled_data = 16'b1101110010110101;
				18'b010000111000010010: oled_data = 16'b1110010011010110;
				18'b010000111010010010: oled_data = 16'b1101010001110100;
				18'b010000111100010010: oled_data = 16'b1101110011010101;
				18'b010000111110010010: oled_data = 16'b1101110011010101;
				18'b010001000000010010: oled_data = 16'b1101110011010101;
				18'b010001000010010010: oled_data = 16'b1101110011010101;
				18'b010001000100010010: oled_data = 16'b1101010001110100;
				18'b010001000110010010: oled_data = 16'b1101110011010101;
				18'b010001001000010010: oled_data = 16'b1101110011010101;
				18'b010001001010010010: oled_data = 16'b1110010011010110;
				18'b010001001100010010: oled_data = 16'b1101010010010101;
				18'b010001001110010010: oled_data = 16'b1100110001010011;
				18'b010001010000010010: oled_data = 16'b1110010011010110;
				18'b010001010010010010: oled_data = 16'b1101110011010101;
				18'b010001010100010010: oled_data = 16'b1101110011010101;
				18'b010001010110010010: oled_data = 16'b1101110011010101;
				18'b010001011000010010: oled_data = 16'b1101110011010101;
				18'b010001011010010010: oled_data = 16'b1110010011110110;
				18'b010001011100010010: oled_data = 16'b1110110101010111;
				18'b010001011110010010: oled_data = 16'b1101110011010101;
				18'b010001100000010010: oled_data = 16'b1101110011010101;
				18'b010001100010010010: oled_data = 16'b1101110011010101;
				18'b010001100100010010: oled_data = 16'b1101110011010110;
				18'b010001100110010010: oled_data = 16'b1101110010110101;
				18'b010001101000010010: oled_data = 16'b1101010010010100;
				18'b010001101010010010: oled_data = 16'b1101010010110100;
				18'b010001101100010010: oled_data = 16'b1110011001011001;
				18'b010001101110010010: oled_data = 16'b1110011001111001;
				18'b010001110000010010: oled_data = 16'b1101010011110101;
				18'b010001110010010010: oled_data = 16'b1101110011010101;
				18'b010001110100010010: oled_data = 16'b1101110011010110;
				18'b010001110110010010: oled_data = 16'b1101010001110100;
				18'b010001111000010010: oled_data = 16'b1011001110010000;
				18'b010001111010010010: oled_data = 16'b1011001110010001;
				18'b010001111100010010: oled_data = 16'b1011101110010001;
				18'b010001111110010010: oled_data = 16'b1101110010110101;
				18'b010010000000010010: oled_data = 16'b1101110011010110;
				18'b010010000010010010: oled_data = 16'b1101110011010110;
				18'b010010000100010010: oled_data = 16'b1101010001110100;
				18'b010010000110010010: oled_data = 16'b1101110011010110;
				18'b010010001000010010: oled_data = 16'b1101110010110101;
				18'b010010001010010010: oled_data = 16'b1101010001110100;
				18'b010010001100010010: oled_data = 16'b1101010001110011;
				18'b010010001110010010: oled_data = 16'b1110010100010100;
				18'b010010010000010010: oled_data = 16'b1101110000110000;
				18'b010010010010010010: oled_data = 16'b1011001001101010;
				18'b010010010100010010: oled_data = 16'b1011001001001001;
				18'b010010010110010010: oled_data = 16'b1011001001001001;
				18'b010010011000010010: oled_data = 16'b1011001001001001;
				18'b010010011010010010: oled_data = 16'b1011001000101001;
				18'b010010011100010010: oled_data = 16'b1011001001001001;
				18'b010010011110010010: oled_data = 16'b1011001000101001;
				18'b010010100000010010: oled_data = 16'b1011001000101001;
				18'b010010100010010010: oled_data = 16'b1011001000101000;
				18'b010010100100010010: oled_data = 16'b1011001000101000;
				18'b010010100110010010: oled_data = 16'b1011001000001000;
				18'b010000011000010011: oled_data = 16'b0101110001110011;
				18'b010000011010010011: oled_data = 16'b0111011000011010;
				18'b010000011100010011: oled_data = 16'b0110110111011001;
				18'b010000011110010011: oled_data = 16'b0111010111111001;
				18'b010000100000010011: oled_data = 16'b1001111011011101;
				18'b010000100010010011: oled_data = 16'b1001111011011100;
				18'b010000100100010011: oled_data = 16'b1000011000111010;
				18'b010000100110010011: oled_data = 16'b0111011001011010;
				18'b010000101000010011: oled_data = 16'b1001010110111001;
				18'b010000101010010011: oled_data = 16'b1101110011010110;
				18'b010000101100010011: oled_data = 16'b1101110011010101;
				18'b010000101110010011: oled_data = 16'b1101110011010101;
				18'b010000110000010011: oled_data = 16'b1101110011010110;
				18'b010000110010010011: oled_data = 16'b1101110011010110;
				18'b010000110100010011: oled_data = 16'b1101010001110100;
				18'b010000110110010011: oled_data = 16'b1101110010110101;
				18'b010000111000010011: oled_data = 16'b1101110011010110;
				18'b010000111010010011: oled_data = 16'b1101010001110100;
				18'b010000111100010011: oled_data = 16'b1101110011010101;
				18'b010000111110010011: oled_data = 16'b1101110011010101;
				18'b010001000000010011: oled_data = 16'b1101110011010101;
				18'b010001000010010011: oled_data = 16'b1101110011010110;
				18'b010001000100010011: oled_data = 16'b1101010001110100;
				18'b010001000110010011: oled_data = 16'b1101110010110101;
				18'b010001001000010011: oled_data = 16'b1101110011010101;
				18'b010001001010010011: oled_data = 16'b1101110011010101;
				18'b010001001100010011: oled_data = 16'b1101110011010101;
				18'b010001001110010011: oled_data = 16'b1100010000010010;
				18'b010001010000010011: oled_data = 16'b1101110011010101;
				18'b010001010010010011: oled_data = 16'b1101110011010101;
				18'b010001010100010011: oled_data = 16'b1101110011010101;
				18'b010001010110010011: oled_data = 16'b1101110011010101;
				18'b010001011000010011: oled_data = 16'b1101110011010101;
				18'b010001011010010011: oled_data = 16'b1101110010110101;
				18'b010001011100010011: oled_data = 16'b1110010011110110;
				18'b010001011110010011: oled_data = 16'b1110010011010110;
				18'b010001100000010011: oled_data = 16'b1101110011010101;
				18'b010001100010010011: oled_data = 16'b1101110011010101;
				18'b010001100100010011: oled_data = 16'b1101110011010101;
				18'b010001100110010011: oled_data = 16'b1101110011010101;
				18'b010001101000010011: oled_data = 16'b1101010001110100;
				18'b010001101010010011: oled_data = 16'b1101110010010100;
				18'b010001101100010011: oled_data = 16'b1101110110110111;
				18'b010001101110010011: oled_data = 16'b1110111100111100;
				18'b010001110000010011: oled_data = 16'b1101111000011000;
				18'b010001110010010011: oled_data = 16'b1101110010110101;
				18'b010001110100010011: oled_data = 16'b1101110011010110;
				18'b010001110110010011: oled_data = 16'b1101110010110101;
				18'b010001111000010011: oled_data = 16'b1101010010110101;
				18'b010001111010010011: oled_data = 16'b1011001111010001;
				18'b010001111100010011: oled_data = 16'b1011001101010000;
				18'b010001111110010011: oled_data = 16'b1011101110110001;
				18'b010010000000010011: oled_data = 16'b1101110011010110;
				18'b010010000010010011: oled_data = 16'b1101110011010110;
				18'b010010000100010011: oled_data = 16'b1101110010010101;
				18'b010010000110010011: oled_data = 16'b1101110010110101;
				18'b010010001000010011: oled_data = 16'b1101010010010100;
				18'b010010001010010011: oled_data = 16'b1100110000110010;
				18'b010010001100010011: oled_data = 16'b1110010100010100;
				18'b010010001110010011: oled_data = 16'b1101110001010001;
				18'b010010010000010011: oled_data = 16'b1011001010001010;
				18'b010010010010010011: oled_data = 16'b1011001001001001;
				18'b010010010100010011: oled_data = 16'b1011001001001001;
				18'b010010010110010011: oled_data = 16'b1011001001001001;
				18'b010010011000010011: oled_data = 16'b1011001001001001;
				18'b010010011010010011: oled_data = 16'b1011001000101001;
				18'b010010011100010011: oled_data = 16'b1011001001001001;
				18'b010010011110010011: oled_data = 16'b1011001000101001;
				18'b010010100000010011: oled_data = 16'b1011001000101001;
				18'b010010100010010011: oled_data = 16'b1011001000101001;
				18'b010010100100010011: oled_data = 16'b1011001000101000;
				18'b010010100110010011: oled_data = 16'b1011001000001000;
				18'b010000011000010100: oled_data = 16'b0110010100010101;
				18'b010000011010010100: oled_data = 16'b0110110111111001;
				18'b010000011100010100: oled_data = 16'b0100110010110101;
				18'b010000011110010100: oled_data = 16'b1000111001011010;
				18'b010000100000010100: oled_data = 16'b1011111101011101;
				18'b010000100010010100: oled_data = 16'b1001011000011010;
				18'b010000100100010100: oled_data = 16'b0101010011010101;
				18'b010000100110010100: oled_data = 16'b0111011000011010;
				18'b010000101000010100: oled_data = 16'b1000011000111010;
				18'b010000101010010100: oled_data = 16'b1101010011010110;
				18'b010000101100010100: oled_data = 16'b1110010011010101;
				18'b010000101110010100: oled_data = 16'b1101110011010110;
				18'b010000110000010100: oled_data = 16'b1101110011010110;
				18'b010000110010010100: oled_data = 16'b1101110011010110;
				18'b010000110100010100: oled_data = 16'b1101010001110100;
				18'b010000110110010100: oled_data = 16'b1101110010110101;
				18'b010000111000010100: oled_data = 16'b1101110011010110;
				18'b010000111010010100: oled_data = 16'b1101010001110100;
				18'b010000111100010100: oled_data = 16'b1101110011010101;
				18'b010000111110010100: oled_data = 16'b1101110011010101;
				18'b010001000000010100: oled_data = 16'b1101110011010101;
				18'b010001000010010100: oled_data = 16'b1101110011010101;
				18'b010001000100010100: oled_data = 16'b1101110010110101;
				18'b010001000110010100: oled_data = 16'b1101110010110101;
				18'b010001001000010100: oled_data = 16'b1101110011010101;
				18'b010001001010010100: oled_data = 16'b1101110011010101;
				18'b010001001100010100: oled_data = 16'b1101110011010101;
				18'b010001001110010100: oled_data = 16'b1100110001110100;
				18'b010001010000010100: oled_data = 16'b1101010010010100;
				18'b010001010010010100: oled_data = 16'b1101110011010110;
				18'b010001010100010100: oled_data = 16'b1101110011010101;
				18'b010001010110010100: oled_data = 16'b1101110011010101;
				18'b010001011000010100: oled_data = 16'b1101110011010101;
				18'b010001011010010100: oled_data = 16'b1101110011010101;
				18'b010001011100010100: oled_data = 16'b1101110011010101;
				18'b010001011110010100: oled_data = 16'b1101110011010110;
				18'b010001100000010100: oled_data = 16'b1101110011010101;
				18'b010001100010010100: oled_data = 16'b1101110011010101;
				18'b010001100100010100: oled_data = 16'b1101110011010101;
				18'b010001100110010100: oled_data = 16'b1101110011010110;
				18'b010001101000010100: oled_data = 16'b1101110010010101;
				18'b010001101010010100: oled_data = 16'b1101010001110100;
				18'b010001101100010100: oled_data = 16'b1101010100010101;
				18'b010001101110010100: oled_data = 16'b1110111011111011;
				18'b010001110000010100: oled_data = 16'b1110111100011011;
				18'b010001110010010100: oled_data = 16'b1101010100110110;
				18'b010001110100010100: oled_data = 16'b1101110010110101;
				18'b010001110110010100: oled_data = 16'b1101110010110101;
				18'b010001111000010100: oled_data = 16'b1101110100010110;
				18'b010001111010010100: oled_data = 16'b1101010101010110;
				18'b010001111100010100: oled_data = 16'b1011001101110000;
				18'b010001111110010100: oled_data = 16'b1011001100110000;
				18'b010010000000010100: oled_data = 16'b1100110000010011;
				18'b010010000010010100: oled_data = 16'b1110010011010110;
				18'b010010000100010100: oled_data = 16'b1101110010010101;
				18'b010010000110010100: oled_data = 16'b1101010010010100;
				18'b010010001000010100: oled_data = 16'b1101010001110011;
				18'b010010001010010100: oled_data = 16'b1101110011010011;
				18'b010010001100010100: oled_data = 16'b1110010011010011;
				18'b010010001110010100: oled_data = 16'b1011101010101011;
				18'b010010010000010100: oled_data = 16'b1011001001001001;
				18'b010010010010010100: oled_data = 16'b1011001001001001;
				18'b010010010100010100: oled_data = 16'b1011001001001001;
				18'b010010010110010100: oled_data = 16'b1011001001001001;
				18'b010010011000010100: oled_data = 16'b1011001001001001;
				18'b010010011010010100: oled_data = 16'b1011001000101001;
				18'b010010011100010100: oled_data = 16'b1011001001001001;
				18'b010010011110010100: oled_data = 16'b1011001000101001;
				18'b010010100000010100: oled_data = 16'b1010101000001000;
				18'b010010100010010100: oled_data = 16'b1011001000101001;
				18'b010010100100010100: oled_data = 16'b1011001000101000;
				18'b010010100110010100: oled_data = 16'b1011001000001000;
				18'b010000011000010101: oled_data = 16'b0110110110010111;
				18'b010000011010010101: oled_data = 16'b0101110101111000;
				18'b010000011100010101: oled_data = 16'b0100010001110101;
				18'b010000011110010101: oled_data = 16'b1001111010011010;
				18'b010000100000010101: oled_data = 16'b1001111010111011;
				18'b010000100010010101: oled_data = 16'b0101010010110110;
				18'b010000100100010101: oled_data = 16'b0100010001010101;
				18'b010000100110010101: oled_data = 16'b0101110101011000;
				18'b010000101000010101: oled_data = 16'b1000011000011001;
				18'b010000101010010101: oled_data = 16'b1101010011010110;
				18'b010000101100010101: oled_data = 16'b1101110011010110;
				18'b010000101110010101: oled_data = 16'b1101110011010101;
				18'b010000110000010101: oled_data = 16'b1101110011010101;
				18'b010000110010010101: oled_data = 16'b1101110011010110;
				18'b010000110100010101: oled_data = 16'b1101010001110100;
				18'b010000110110010101: oled_data = 16'b1101110010110101;
				18'b010000111000010101: oled_data = 16'b1101110011010101;
				18'b010000111010010101: oled_data = 16'b1100110000110011;
				18'b010000111100010101: oled_data = 16'b1101110011010101;
				18'b010000111110010101: oled_data = 16'b1101110011010101;
				18'b010001000000010101: oled_data = 16'b1101110011010101;
				18'b010001000010010101: oled_data = 16'b1101110011010101;
				18'b010001000100010101: oled_data = 16'b1101110010110101;
				18'b010001000110010101: oled_data = 16'b1101010010010100;
				18'b010001001000010101: oled_data = 16'b1101110011010110;
				18'b010001001010010101: oled_data = 16'b1101110011010101;
				18'b010001001100010101: oled_data = 16'b1101110011010101;
				18'b010001001110010101: oled_data = 16'b1101010010110101;
				18'b010001010000010101: oled_data = 16'b1100110001110100;
				18'b010001010010010101: oled_data = 16'b1101110011010110;
				18'b010001010100010101: oled_data = 16'b1101110011010101;
				18'b010001010110010101: oled_data = 16'b1101110011010101;
				18'b010001011000010101: oled_data = 16'b1101110011010101;
				18'b010001011010010101: oled_data = 16'b1101110011010101;
				18'b010001011100010101: oled_data = 16'b1101110011010101;
				18'b010001011110010101: oled_data = 16'b1101110011010101;
				18'b010001100000010101: oled_data = 16'b1110010011010110;
				18'b010001100010010101: oled_data = 16'b1110010011010110;
				18'b010001100100010101: oled_data = 16'b1101110011010101;
				18'b010001100110010101: oled_data = 16'b1101110011010101;
				18'b010001101000010101: oled_data = 16'b1101110011010101;
				18'b010001101010010101: oled_data = 16'b1101010001110100;
				18'b010001101100010101: oled_data = 16'b1101010010010100;
				18'b010001101110010101: oled_data = 16'b1101111010011010;
				18'b010001110000010101: oled_data = 16'b1101111011011010;
				18'b010001110010010101: oled_data = 16'b1101011000111000;
				18'b010001110100010101: oled_data = 16'b1101010011110110;
				18'b010001110110010101: oled_data = 16'b1101110011010101;
				18'b010001111000010101: oled_data = 16'b1101010011010101;
				18'b010001111010010101: oled_data = 16'b1101110111111000;
				18'b010001111100010101: oled_data = 16'b1011001110010000;
				18'b010001111110010101: oled_data = 16'b1011001101010000;
				18'b010010000000010101: oled_data = 16'b1011001110010001;
				18'b010010000010010101: oled_data = 16'b1101110010010101;
				18'b010010000100010101: oled_data = 16'b1101110010110101;
				18'b010010000110010101: oled_data = 16'b1011101110110001;
				18'b010010001000010101: oled_data = 16'b1101110010110011;
				18'b010010001010010101: oled_data = 16'b1110110100010100;
				18'b010010001100010101: oled_data = 16'b1100001100101101;
				18'b010010001110010101: oled_data = 16'b1011001000101001;
				18'b010010010000010101: oled_data = 16'b1011101001001001;
				18'b010010010010010101: oled_data = 16'b1011101000101001;
				18'b010010010100010101: oled_data = 16'b1011001001001001;
				18'b010010010110010101: oled_data = 16'b1011001001001001;
				18'b010010011000010101: oled_data = 16'b1011001001001001;
				18'b010010011010010101: oled_data = 16'b1011001001001001;
				18'b010010011100010101: oled_data = 16'b1011001000101001;
				18'b010010011110010101: oled_data = 16'b1010001000001000;
				18'b010010100000010101: oled_data = 16'b1010101000001000;
				18'b010010100010010101: oled_data = 16'b1011001000101001;
				18'b010010100100010101: oled_data = 16'b1011001000101000;
				18'b010010100110010101: oled_data = 16'b1011001000001000;
				18'b010000011000010110: oled_data = 16'b0111010111111001;
				18'b010000011010010110: oled_data = 16'b0101010100010111;
				18'b010000011100010110: oled_data = 16'b0100110001010101;
				18'b010000011110010110: oled_data = 16'b1001011001111011;
				18'b010000100000010110: oled_data = 16'b0110110100110111;
				18'b010000100010010110: oled_data = 16'b0100010001010101;
				18'b010000100100010110: oled_data = 16'b0100010001110110;
				18'b010000100110010110: oled_data = 16'b0100110011010110;
				18'b010000101000010110: oled_data = 16'b1000010111111001;
				18'b010000101010010110: oled_data = 16'b1101010011010110;
				18'b010000101100010110: oled_data = 16'b1101110011010101;
				18'b010000101110010110: oled_data = 16'b1101110011010101;
				18'b010000110000010110: oled_data = 16'b1101110011010101;
				18'b010000110010010110: oled_data = 16'b1101110011010110;
				18'b010000110100010110: oled_data = 16'b1101010001110100;
				18'b010000110110010110: oled_data = 16'b1101110010110101;
				18'b010000111000010110: oled_data = 16'b1101110011010101;
				18'b010000111010010110: oled_data = 16'b1100110000010011;
				18'b010000111100010110: oled_data = 16'b1101110011010101;
				18'b010000111110010110: oled_data = 16'b1101110011010101;
				18'b010001000000010110: oled_data = 16'b1101110011010101;
				18'b010001000010010110: oled_data = 16'b1101110011010101;
				18'b010001000100010110: oled_data = 16'b1101110011010110;
				18'b010001000110010110: oled_data = 16'b1100110001010011;
				18'b010001001000010110: oled_data = 16'b1101110011010101;
				18'b010001001010010110: oled_data = 16'b1101110011010101;
				18'b010001001100010110: oled_data = 16'b1101110011010101;
				18'b010001001110010110: oled_data = 16'b1101110011010101;
				18'b010001010000010110: oled_data = 16'b1101010010010100;
				18'b010001010010010110: oled_data = 16'b1101010010110101;
				18'b010001010100010110: oled_data = 16'b1101110011010101;
				18'b010001010110010110: oled_data = 16'b1101110011010101;
				18'b010001011000010110: oled_data = 16'b1101110011010101;
				18'b010001011010010110: oled_data = 16'b1101110011010101;
				18'b010001011100010110: oled_data = 16'b1110010011010101;
				18'b010001011110010110: oled_data = 16'b1110010011010101;
				18'b010001100000010110: oled_data = 16'b1110010011010110;
				18'b010001100010010110: oled_data = 16'b1110010011010110;
				18'b010001100100010110: oled_data = 16'b1110010011010110;
				18'b010001100110010110: oled_data = 16'b1110010011010110;
				18'b010001101000010110: oled_data = 16'b1110010011010110;
				18'b010001101010010110: oled_data = 16'b1101010010010101;
				18'b010001101100010110: oled_data = 16'b1100110001010100;
				18'b010001101110010110: oled_data = 16'b1100110111010111;
				18'b010001110000010110: oled_data = 16'b1101011010011001;
				18'b010001110010010110: oled_data = 16'b1110111101011100;
				18'b010001110100010110: oled_data = 16'b1010110010110011;
				18'b010001110110010110: oled_data = 16'b1101010010110101;
				18'b010001111000010110: oled_data = 16'b1101110011010101;
				18'b010001111010010110: oled_data = 16'b1101010110110111;
				18'b010001111100010110: oled_data = 16'b1100010001010011;
				18'b010001111110010110: oled_data = 16'b1010101100001111;
				18'b010010000000010110: oled_data = 16'b1011001101110000;
				18'b010010000010010110: oled_data = 16'b1100001111110010;
				18'b010010000100010110: oled_data = 16'b1101110010110101;
				18'b010010000110010110: oled_data = 16'b1100010000010010;
				18'b010010001000010110: oled_data = 16'b1110110100010100;
				18'b010010001010010110: oled_data = 16'b1101010000001111;
				18'b010010001100010110: oled_data = 16'b1011001001001001;
				18'b010010001110010110: oled_data = 16'b1011101001001001;
				18'b010010010000010110: oled_data = 16'b1011101001001001;
				18'b010010010010010110: oled_data = 16'b1011101001001001;
				18'b010010010100010110: oled_data = 16'b1011001001001001;
				18'b010010010110010110: oled_data = 16'b1011001001001001;
				18'b010010011000010110: oled_data = 16'b1011001001001001;
				18'b010010011010010110: oled_data = 16'b1010101000101000;
				18'b010010011100010110: oled_data = 16'b1010001000001000;
				18'b010010011110010110: oled_data = 16'b1011001000101001;
				18'b010010100000010110: oled_data = 16'b1011001000101001;
				18'b010010100010010110: oled_data = 16'b1011001000101001;
				18'b010010100100010110: oled_data = 16'b1011001000101000;
				18'b010010100110010110: oled_data = 16'b1011001000001000;
				18'b010000011000010111: oled_data = 16'b0111011000011010;
				18'b010000011010010111: oled_data = 16'b0101010011010110;
				18'b010000011100010111: oled_data = 16'b0100110001010101;
				18'b010000011110010111: oled_data = 16'b0110010100011000;
				18'b010000100000010111: oled_data = 16'b0101010001110110;
				18'b010000100010010111: oled_data = 16'b0100110001010110;
				18'b010000100100010111: oled_data = 16'b0100010001110101;
				18'b010000100110010111: oled_data = 16'b0100110010110110;
				18'b010000101000010111: oled_data = 16'b1000110110011001;
				18'b010000101010010111: oled_data = 16'b1101110011010110;
				18'b010000101100010111: oled_data = 16'b1101110011010101;
				18'b010000101110010111: oled_data = 16'b1101110011010101;
				18'b010000110000010111: oled_data = 16'b1101110011010101;
				18'b010000110010010111: oled_data = 16'b1101110011010110;
				18'b010000110100010111: oled_data = 16'b1101010010010100;
				18'b010000110110010111: oled_data = 16'b1101110010110101;
				18'b010000111000010111: oled_data = 16'b1101110011010101;
				18'b010000111010010111: oled_data = 16'b1100110000010011;
				18'b010000111100010111: oled_data = 16'b1101110011010101;
				18'b010000111110010111: oled_data = 16'b1101110011010101;
				18'b010001000000010111: oled_data = 16'b1101110011010101;
				18'b010001000010010111: oled_data = 16'b1101110011010101;
				18'b010001000100010111: oled_data = 16'b1101110011010110;
				18'b010001000110010111: oled_data = 16'b1100110001110100;
				18'b010001001000010111: oled_data = 16'b1101010010010101;
				18'b010001001010010111: oled_data = 16'b1101110011010110;
				18'b010001001100010111: oled_data = 16'b1101110011010101;
				18'b010001001110010111: oled_data = 16'b1101110011010101;
				18'b010001010000010111: oled_data = 16'b1101010010110101;
				18'b010001010010010111: oled_data = 16'b1100110010110100;
				18'b010001010100010111: oled_data = 16'b1101110011010101;
				18'b010001010110010111: oled_data = 16'b1101110011010101;
				18'b010001011000010111: oled_data = 16'b1110010011010101;
				18'b010001011010010111: oled_data = 16'b1101110011010101;
				18'b010001011100010111: oled_data = 16'b1110010011010101;
				18'b010001011110010111: oled_data = 16'b1101110011010101;
				18'b010001100000010111: oled_data = 16'b1101110011010101;
				18'b010001100010010111: oled_data = 16'b1101110011010101;
				18'b010001100100010111: oled_data = 16'b1101110011010101;
				18'b010001100110010111: oled_data = 16'b1101110010110101;
				18'b010001101000010111: oled_data = 16'b1101010010010100;
				18'b010001101010010111: oled_data = 16'b1101010001110100;
				18'b010001101100010111: oled_data = 16'b1100110000110011;
				18'b010001101110010111: oled_data = 16'b1101010101110110;
				18'b010001110000010111: oled_data = 16'b1111011101111100;
				18'b010001110010010111: oled_data = 16'b1101011001111001;
				18'b010001110100010111: oled_data = 16'b0110101011101011;
				18'b010001110110010111: oled_data = 16'b1100110011010100;
				18'b010001111000010111: oled_data = 16'b1101110011010110;
				18'b010001111010010111: oled_data = 16'b1101010101010111;
				18'b010001111100010111: oled_data = 16'b1100110011010101;
				18'b010001111110010111: oled_data = 16'b1011001100110000;
				18'b010010000000010111: oled_data = 16'b1011001101010000;
				18'b010010000010010111: oled_data = 16'b1011101110010001;
				18'b010010000100010111: oled_data = 16'b1100110000110010;
				18'b010010000110010111: oled_data = 16'b1110010011110100;
				18'b010010001000010111: oled_data = 16'b1110010010110010;
				18'b010010001010010111: oled_data = 16'b1011101010001010;
				18'b010010001100010111: oled_data = 16'b1011001001001001;
				18'b010010001110010111: oled_data = 16'b1011001001001001;
				18'b010010010000010111: oled_data = 16'b1011001001001001;
				18'b010010010010010111: oled_data = 16'b1011001001001001;
				18'b010010010100010111: oled_data = 16'b1011001001001001;
				18'b010010010110010111: oled_data = 16'b1011001001001001;
				18'b010010011000010111: oled_data = 16'b1011001000101001;
				18'b010010011010010111: oled_data = 16'b1010001000001000;
				18'b010010011100010111: oled_data = 16'b1011001001001001;
				18'b010010011110010111: oled_data = 16'b1011001000101001;
				18'b010010100000010111: oled_data = 16'b1011001000101001;
				18'b010010100010010111: oled_data = 16'b1011001000101001;
				18'b010010100100010111: oled_data = 16'b1011001000101000;
				18'b010010100110010111: oled_data = 16'b1011001000001000;
				18'b010000011000011000: oled_data = 16'b0111011000011010;
				18'b010000011010011000: oled_data = 16'b0101010010110110;
				18'b010000011100011000: oled_data = 16'b0100110001010110;
				18'b010000011110011000: oled_data = 16'b0100110001010110;
				18'b010000100000011000: oled_data = 16'b0100110001110110;
				18'b010000100010011000: oled_data = 16'b0100110001010110;
				18'b010000100100011000: oled_data = 16'b0100110001010101;
				18'b010000100110011000: oled_data = 16'b0101010011010110;
				18'b010000101000011000: oled_data = 16'b1001110100111000;
				18'b010000101010011000: oled_data = 16'b1101110010110110;
				18'b010000101100011000: oled_data = 16'b1101110011010101;
				18'b010000101110011000: oled_data = 16'b1101110011010101;
				18'b010000110000011000: oled_data = 16'b1101110011010101;
				18'b010000110010011000: oled_data = 16'b1101110011010110;
				18'b010000110100011000: oled_data = 16'b1101010010010100;
				18'b010000110110011000: oled_data = 16'b1101110010110101;
				18'b010000111000011000: oled_data = 16'b1101110011010101;
				18'b010000111010011000: oled_data = 16'b1100110000110011;
				18'b010000111100011000: oled_data = 16'b1101110010110101;
				18'b010000111110011000: oled_data = 16'b1101110011010101;
				18'b010001000000011000: oled_data = 16'b1101110011010101;
				18'b010001000010011000: oled_data = 16'b1101110011010101;
				18'b010001000100011000: oled_data = 16'b1101110011010110;
				18'b010001000110011000: oled_data = 16'b1101010010110101;
				18'b010001001000011000: oled_data = 16'b1100110001110100;
				18'b010001001010011000: oled_data = 16'b1101110011010101;
				18'b010001001100011000: oled_data = 16'b1101110011010101;
				18'b010001001110011000: oled_data = 16'b1101110011010101;
				18'b010001010000011000: oled_data = 16'b1101110010110101;
				18'b010001010010011000: oled_data = 16'b1101010101110110;
				18'b010001010100011000: oled_data = 16'b1101010011010101;
				18'b010001010110011000: oled_data = 16'b1110010011010101;
				18'b010001011000011000: oled_data = 16'b1110010011010101;
				18'b010001011010011000: oled_data = 16'b1101110011010101;
				18'b010001011100011000: oled_data = 16'b1110010011010101;
				18'b010001011110011000: oled_data = 16'b1101110011010101;
				18'b010001100000011000: oled_data = 16'b1101110011010101;
				18'b010001100010011000: oled_data = 16'b1101110011010101;
				18'b010001100100011000: oled_data = 16'b1101110011010101;
				18'b010001100110011000: oled_data = 16'b1101110010110101;
				18'b010001101000011000: oled_data = 16'b1101110010110101;
				18'b010001101010011000: oled_data = 16'b1101110011010101;
				18'b010001101100011000: oled_data = 16'b1101010010010100;
				18'b010001101110011000: oled_data = 16'b1100110101010110;
				18'b010001110000011000: oled_data = 16'b1110111101011100;
				18'b010001110010011000: oled_data = 16'b1001010010010001;
				18'b010001110100011000: oled_data = 16'b0100000111000110;
				18'b010001110110011000: oled_data = 16'b1011110110010110;
				18'b010001111000011000: oled_data = 16'b1101110100110110;
				18'b010001111010011000: oled_data = 16'b1101110100110110;
				18'b010001111100011000: oled_data = 16'b1101010101010111;
				18'b010001111110011000: oled_data = 16'b1011001101110000;
				18'b010010000000011000: oled_data = 16'b1010101100001111;
				18'b010010000010011000: oled_data = 16'b1011001101110001;
				18'b010010000100011000: oled_data = 16'b1101010001110010;
				18'b010010000110011000: oled_data = 16'b1110110100010100;
				18'b010010001000011000: oled_data = 16'b1100101101101101;
				18'b010010001010011000: oled_data = 16'b1011001000101001;
				18'b010010001100011000: oled_data = 16'b1011101001001001;
				18'b010010001110011000: oled_data = 16'b1011001001001001;
				18'b010010010000011000: oled_data = 16'b1011001001001001;
				18'b010010010010011000: oled_data = 16'b1011001001001001;
				18'b010010010100011000: oled_data = 16'b1011001001001001;
				18'b010010010110011000: oled_data = 16'b1011001000101001;
				18'b010010011000011000: oled_data = 16'b1010101000001000;
				18'b010010011010011000: oled_data = 16'b1011001000101001;
				18'b010010011100011000: oled_data = 16'b1011001001001001;
				18'b010010011110011000: oled_data = 16'b1011001000101001;
				18'b010010100000011000: oled_data = 16'b1011001000101001;
				18'b010010100010011000: oled_data = 16'b1011001000101001;
				18'b010010100100011000: oled_data = 16'b1011001000101000;
				18'b010010100110011000: oled_data = 16'b1010101000001000;
				18'b010000011000011001: oled_data = 16'b0111011000111010;
				18'b010000011010011001: oled_data = 16'b0101110100010111;
				18'b010000011100011001: oled_data = 16'b0100010001010101;
				18'b010000011110011001: oled_data = 16'b0100110001010110;
				18'b010000100000011001: oled_data = 16'b0100110001110101;
				18'b010000100010011001: oled_data = 16'b0100110001010101;
				18'b010000100100011001: oled_data = 16'b0100010001010101;
				18'b010000100110011001: oled_data = 16'b0110010100111000;
				18'b010000101000011001: oled_data = 16'b1010110101011000;
				18'b010000101010011001: oled_data = 16'b1110010011010101;
				18'b010000101100011001: oled_data = 16'b1101110011010101;
				18'b010000101110011001: oled_data = 16'b1101110011010101;
				18'b010000110000011001: oled_data = 16'b1101110011010101;
				18'b010000110010011001: oled_data = 16'b1101110011010110;
				18'b010000110100011001: oled_data = 16'b1101010010010101;
				18'b010000110110011001: oled_data = 16'b1101110010110101;
				18'b010000111000011001: oled_data = 16'b1101110011010110;
				18'b010000111010011001: oled_data = 16'b1101010001010100;
				18'b010000111100011001: oled_data = 16'b1101110010110101;
				18'b010000111110011001: oled_data = 16'b1101110011010101;
				18'b010001000000011001: oled_data = 16'b1101110011010101;
				18'b010001000010011001: oled_data = 16'b1101110011010101;
				18'b010001000100011001: oled_data = 16'b1101110011010101;
				18'b010001000110011001: oled_data = 16'b1101110011010101;
				18'b010001001000011001: oled_data = 16'b1101010011110101;
				18'b010001001010011001: oled_data = 16'b1101010010010100;
				18'b010001001100011001: oled_data = 16'b1101110011010101;
				18'b010001001110011001: oled_data = 16'b1101110011010101;
				18'b010001010000011001: oled_data = 16'b1101110011010101;
				18'b010001010010011001: oled_data = 16'b1101010101010110;
				18'b010001010100011001: oled_data = 16'b1110011000011000;
				18'b010001010110011001: oled_data = 16'b1101010010110101;
				18'b010001011000011001: oled_data = 16'b1101110011010101;
				18'b010001011010011001: oled_data = 16'b1101110011010110;
				18'b010001011100011001: oled_data = 16'b1101110011010101;
				18'b010001011110011001: oled_data = 16'b1101110011010101;
				18'b010001100000011001: oled_data = 16'b1101110011010101;
				18'b010001100010011001: oled_data = 16'b1101110011010101;
				18'b010001100100011001: oled_data = 16'b1101110011010101;
				18'b010001100110011001: oled_data = 16'b1101110011010101;
				18'b010001101000011001: oled_data = 16'b1101110011010101;
				18'b010001101010011001: oled_data = 16'b1101110011010110;
				18'b010001101100011001: oled_data = 16'b1101010010010100;
				18'b010001101110011001: oled_data = 16'b1100110100010101;
				18'b010001110000011001: oled_data = 16'b1101111001111001;
				18'b010001110010011001: oled_data = 16'b0101101001101001;
				18'b010001110100011001: oled_data = 16'b0101001001101001;
				18'b010001110110011001: oled_data = 16'b1101111010111010;
				18'b010001111000011001: oled_data = 16'b1101010110110111;
				18'b010001111010011001: oled_data = 16'b1101110011110110;
				18'b010001111100011001: oled_data = 16'b1101110110111000;
				18'b010001111110011001: oled_data = 16'b1011001110010001;
				18'b010010000000011001: oled_data = 16'b1011001101110001;
				18'b010010000010011001: oled_data = 16'b1100001111010001;
				18'b010010000100011001: oled_data = 16'b1110110011110100;
				18'b010010000110011001: oled_data = 16'b1101110001110010;
				18'b010010001000011001: oled_data = 16'b1011101001101010;
				18'b010010001010011001: oled_data = 16'b1011001001001001;
				18'b010010001100011001: oled_data = 16'b1011001001001001;
				18'b010010001110011001: oled_data = 16'b1011001001001001;
				18'b010010010000011001: oled_data = 16'b1011001001001001;
				18'b010010010010011001: oled_data = 16'b1011001001001001;
				18'b010010010100011001: oled_data = 16'b1011001000101001;
				18'b010010010110011001: oled_data = 16'b1010101000001000;
				18'b010010011000011001: oled_data = 16'b1011001000101001;
				18'b010010011010011001: oled_data = 16'b1011001001001001;
				18'b010010011100011001: oled_data = 16'b1011001000101001;
				18'b010010011110011001: oled_data = 16'b1011001000101001;
				18'b010010100000011001: oled_data = 16'b1011001000101001;
				18'b010010100010011001: oled_data = 16'b1011001000101000;
				18'b010010100100011001: oled_data = 16'b1011001000101000;
				18'b010010100110011001: oled_data = 16'b1010101000101000;
				18'b010000011000011010: oled_data = 16'b0111011000111011;
				18'b010000011010011010: oled_data = 16'b0110110110111001;
				18'b010000011100011010: oled_data = 16'b0100010001110101;
				18'b010000011110011010: oled_data = 16'b0100110001010101;
				18'b010000100000011010: oled_data = 16'b0100010001010101;
				18'b010000100010011010: oled_data = 16'b0100010001010101;
				18'b010000100100011010: oled_data = 16'b0100110010010110;
				18'b010000100110011010: oled_data = 16'b0110110111111010;
				18'b010000101000011010: oled_data = 16'b1010010100010111;
				18'b010000101010011010: oled_data = 16'b1110010011010101;
				18'b010000101100011010: oled_data = 16'b1101110011010110;
				18'b010000101110011010: oled_data = 16'b1101110011010101;
				18'b010000110000011010: oled_data = 16'b1101110011010101;
				18'b010000110010011010: oled_data = 16'b1101110011010110;
				18'b010000110100011010: oled_data = 16'b1101110010010101;
				18'b010000110110011010: oled_data = 16'b1101110010110101;
				18'b010000111000011010: oled_data = 16'b1101110011010110;
				18'b010000111010011010: oled_data = 16'b1100110001010011;
				18'b010000111100011010: oled_data = 16'b1101010010010101;
				18'b010000111110011010: oled_data = 16'b1101110011010110;
				18'b010001000000011010: oled_data = 16'b1101110011010101;
				18'b010001000010011010: oled_data = 16'b1101110011010101;
				18'b010001000100011010: oled_data = 16'b1101110011010101;
				18'b010001000110011010: oled_data = 16'b1101110011010101;
				18'b010001001000011010: oled_data = 16'b1101110111011000;
				18'b010001001010011010: oled_data = 16'b1101010100110110;
				18'b010001001100011010: oled_data = 16'b1101110010110101;
				18'b010001001110011010: oled_data = 16'b1101110011010101;
				18'b010001010000011010: oled_data = 16'b1101110011010101;
				18'b010001010010011010: oled_data = 16'b1101010011010101;
				18'b010001010100011010: oled_data = 16'b1110111001011010;
				18'b010001010110011010: oled_data = 16'b1101110110110111;
				18'b010001011000011010: oled_data = 16'b1101010010110101;
				18'b010001011010011010: oled_data = 16'b1101110010010101;
				18'b010001011100011010: oled_data = 16'b1101110011010110;
				18'b010001011110011010: oled_data = 16'b1101110011010101;
				18'b010001100000011010: oled_data = 16'b1101110011010101;
				18'b010001100010011010: oled_data = 16'b1101110011010101;
				18'b010001100100011010: oled_data = 16'b1101110011010101;
				18'b010001100110011010: oled_data = 16'b1101110011010101;
				18'b010001101000011010: oled_data = 16'b1101110011010101;
				18'b010001101010011010: oled_data = 16'b1101110011010110;
				18'b010001101100011010: oled_data = 16'b1101110010010101;
				18'b010001101110011010: oled_data = 16'b1100110011110100;
				18'b010001110000011010: oled_data = 16'b1010110011010011;
				18'b010001110010011010: oled_data = 16'b0011100110000110;
				18'b010001110100011010: oled_data = 16'b1001110010010010;
				18'b010001110110011010: oled_data = 16'b1110011100011011;
				18'b010001111000011010: oled_data = 16'b1101111010011010;
				18'b010001111010011010: oled_data = 16'b1101010100110110;
				18'b010001111100011010: oled_data = 16'b1110011001111010;
				18'b010001111110011010: oled_data = 16'b1011001111110010;
				18'b010010000000011010: oled_data = 16'b1011001110010000;
				18'b010010000010011010: oled_data = 16'b1101110010110011;
				18'b010010000100011010: oled_data = 16'b1110110100010100;
				18'b010010000110011010: oled_data = 16'b1100101100101101;
				18'b010010001000011010: oled_data = 16'b1011001001001001;
				18'b010010001010011010: oled_data = 16'b1011001001001001;
				18'b010010001100011010: oled_data = 16'b1011001001001001;
				18'b010010001110011010: oled_data = 16'b1011001001001001;
				18'b010010010000011010: oled_data = 16'b1011001001001001;
				18'b010010010010011010: oled_data = 16'b1011001001001001;
				18'b010010010100011010: oled_data = 16'b1010101000001000;
				18'b010010010110011010: oled_data = 16'b1011001000101001;
				18'b010010011000011010: oled_data = 16'b1011001001001001;
				18'b010010011010011010: oled_data = 16'b1011001001001001;
				18'b010010011100011010: oled_data = 16'b1011001000101001;
				18'b010010011110011010: oled_data = 16'b1011001000101001;
				18'b010010100000011010: oled_data = 16'b1011001000101001;
				18'b010010100010011010: oled_data = 16'b1011001000101000;
				18'b010010100100011010: oled_data = 16'b1011001000101000;
				18'b010010100110011010: oled_data = 16'b1010101000101000;
				18'b010000011000011011: oled_data = 16'b0110110110110111;
				18'b010000011010011011: oled_data = 16'b0111011000011001;
				18'b010000011100011011: oled_data = 16'b0101110101010111;
				18'b010000011110011011: oled_data = 16'b0100110001110101;
				18'b010000100000011011: oled_data = 16'b0100110001110101;
				18'b010000100010011011: oled_data = 16'b0100110010110110;
				18'b010000100100011011: oled_data = 16'b0110110110111010;
				18'b010000100110011011: oled_data = 16'b0111011000111010;
				18'b010000101000011011: oled_data = 16'b1011010010110101;
				18'b010000101010011011: oled_data = 16'b1101110010010101;
				18'b010000101100011011: oled_data = 16'b1101010001110100;
				18'b010000101110011011: oled_data = 16'b1101010010010101;
				18'b010000110000011011: oled_data = 16'b1101110010110101;
				18'b010000110010011011: oled_data = 16'b1110010011010110;
				18'b010000110100011011: oled_data = 16'b1101110010010101;
				18'b010000110110011011: oled_data = 16'b1101110010010101;
				18'b010000111000011011: oled_data = 16'b1110010011010110;
				18'b010000111010011011: oled_data = 16'b1101010001110100;
				18'b010000111100011011: oled_data = 16'b1101010010010100;
				18'b010000111110011011: oled_data = 16'b1101110011010110;
				18'b010001000000011011: oled_data = 16'b1101110011010101;
				18'b010001000010011011: oled_data = 16'b1101110011010101;
				18'b010001000100011011: oled_data = 16'b1101110011010101;
				18'b010001000110011011: oled_data = 16'b1101110010110101;
				18'b010001001000011011: oled_data = 16'b1101110111010111;
				18'b010001001010011011: oled_data = 16'b1110111010111010;
				18'b010001001100011011: oled_data = 16'b1100110011110101;
				18'b010001001110011011: oled_data = 16'b1101110010110101;
				18'b010001010000011011: oled_data = 16'b1101110011010110;
				18'b010001010010011011: oled_data = 16'b1101110010110101;
				18'b010001010100011011: oled_data = 16'b1101110101110111;
				18'b010001010110011011: oled_data = 16'b1110111011011011;
				18'b010001011000011011: oled_data = 16'b1100110100010101;
				18'b010001011010011011: oled_data = 16'b1101010001110100;
				18'b010001011100011011: oled_data = 16'b1110010011010110;
				18'b010001011110011011: oled_data = 16'b1101110011010101;
				18'b010001100000011011: oled_data = 16'b1101110011010101;
				18'b010001100010011011: oled_data = 16'b1101110011010101;
				18'b010001100100011011: oled_data = 16'b1101110011010101;
				18'b010001100110011011: oled_data = 16'b1101110011010101;
				18'b010001101000011011: oled_data = 16'b1101110011010101;
				18'b010001101010011011: oled_data = 16'b1101110011010101;
				18'b010001101100011011: oled_data = 16'b1101110010110101;
				18'b010001101110011011: oled_data = 16'b1100110010010011;
				18'b010001110000011011: oled_data = 16'b0110001011001010;
				18'b010001110010011011: oled_data = 16'b0100101000001000;
				18'b010001110100011011: oled_data = 16'b1101111010011001;
				18'b010001110110011011: oled_data = 16'b1110011011111011;
				18'b010001111000011011: oled_data = 16'b1110011011111011;
				18'b010001111010011011: oled_data = 16'b1101010111110111;
				18'b010001111100011011: oled_data = 16'b1110011011011010;
				18'b010001111110011011: oled_data = 16'b1100010011110101;
				18'b010010000000011011: oled_data = 16'b1011001110010000;
				18'b010010000010011011: oled_data = 16'b1110010100010100;
				18'b010010000100011011: oled_data = 16'b1101110001110001;
				18'b010010000110011011: oled_data = 16'b1011101001101010;
				18'b010010001000011011: oled_data = 16'b1011101001001001;
				18'b010010001010011011: oled_data = 16'b1100001011001100;
				18'b010010001100011011: oled_data = 16'b1011101001101010;
				18'b010010001110011011: oled_data = 16'b1011001001001001;
				18'b010010010000011011: oled_data = 16'b1011001001001001;
				18'b010010010010011011: oled_data = 16'b1011001000101000;
				18'b010010010100011011: oled_data = 16'b1010101000101001;
				18'b010010010110011011: oled_data = 16'b1011001001001001;
				18'b010010011000011011: oled_data = 16'b1011001001001001;
				18'b010010011010011011: oled_data = 16'b1011001000101001;
				18'b010010011100011011: oled_data = 16'b1011001000101001;
				18'b010010011110011011: oled_data = 16'b1011001000101001;
				18'b010010100000011011: oled_data = 16'b1011001000101001;
				18'b010010100010011011: oled_data = 16'b1011001000101000;
				18'b010010100100011011: oled_data = 16'b1011001000101000;
				18'b010010100110011011: oled_data = 16'b1010101000101000;
				18'b010000011000011100: oled_data = 16'b0011001010001100;
				18'b010000011010011100: oled_data = 16'b0101110001110010;
				18'b010000011100011100: oled_data = 16'b0110110111111001;
				18'b010000011110011100: oled_data = 16'b0110110110111010;
				18'b010000100000011100: oled_data = 16'b0110110110111001;
				18'b010000100010011100: oled_data = 16'b0111010111111010;
				18'b010000100100011100: oled_data = 16'b0111111000111011;
				18'b010000100110011100: oled_data = 16'b0111010111111010;
				18'b010000101000011100: oled_data = 16'b1011110010010101;
				18'b010000101010011100: oled_data = 16'b1101110010110101;
				18'b010000101100011100: oled_data = 16'b1101110011010110;
				18'b010000101110011100: oled_data = 16'b1110010011010110;
				18'b010000110000011100: oled_data = 16'b1101010010010100;
				18'b010000110010011100: oled_data = 16'b1101110011010101;
				18'b010000110100011100: oled_data = 16'b1101110010110101;
				18'b010000110110011100: oled_data = 16'b1101110010010101;
				18'b010000111000011100: oled_data = 16'b1110010011010110;
				18'b010000111010011100: oled_data = 16'b1101010010010100;
				18'b010000111100011100: oled_data = 16'b1101010010010101;
				18'b010000111110011100: oled_data = 16'b1101110011010101;
				18'b010001000000011100: oled_data = 16'b1101110011010101;
				18'b010001000010011100: oled_data = 16'b1101110011010101;
				18'b010001000100011100: oled_data = 16'b1101110011010101;
				18'b010001000110011100: oled_data = 16'b1101110011010101;
				18'b010001001000011100: oled_data = 16'b1101010101110110;
				18'b010001001010011100: oled_data = 16'b1110111100011011;
				18'b010001001100011100: oled_data = 16'b1110011001111001;
				18'b010001001110011100: oled_data = 16'b1101010011010101;
				18'b010001010000011100: oled_data = 16'b1101110010110101;
				18'b010001010010011100: oled_data = 16'b1110010010110101;
				18'b010001010100011100: oled_data = 16'b1101110011110101;
				18'b010001010110011100: oled_data = 16'b1110111010011010;
				18'b010001011000011100: oled_data = 16'b1101111000111000;
				18'b010001011010011100: oled_data = 16'b1100110100010101;
				18'b010001011100011100: oled_data = 16'b1101110010110101;
				18'b010001011110011100: oled_data = 16'b1101110011010101;
				18'b010001100000011100: oled_data = 16'b1101110011010101;
				18'b010001100010011100: oled_data = 16'b1101110011010101;
				18'b010001100100011100: oled_data = 16'b1101110011010101;
				18'b010001100110011100: oled_data = 16'b1101110011010101;
				18'b010001101000011100: oled_data = 16'b1101110011010101;
				18'b010001101010011100: oled_data = 16'b1101110011010101;
				18'b010001101100011100: oled_data = 16'b1110010011010110;
				18'b010001101110011100: oled_data = 16'b1010101110110000;
				18'b010001110000011100: oled_data = 16'b0011100101100101;
				18'b010001110010011100: oled_data = 16'b1001010000110000;
				18'b010001110100011100: oled_data = 16'b1110111100111011;
				18'b010001110110011100: oled_data = 16'b1110111100011010;
				18'b010001111000011100: oled_data = 16'b1110111100111011;
				18'b010001111010011100: oled_data = 16'b1110011011111010;
				18'b010001111100011100: oled_data = 16'b1110011011111010;
				18'b010001111110011100: oled_data = 16'b1101010111010111;
				18'b010010000000011100: oled_data = 16'b1100010000110001;
				18'b010010000010011100: oled_data = 16'b1110110100010100;
				18'b010010000100011100: oled_data = 16'b1100101101101101;
				18'b010010000110011100: oled_data = 16'b1011001000101001;
				18'b010010001000011100: oled_data = 16'b1011101010001010;
				18'b010010001010011100: oled_data = 16'b1101001110001110;
				18'b010010001100011100: oled_data = 16'b1011001001001010;
				18'b010010001110011100: oled_data = 16'b1011101001001001;
				18'b010010010000011100: oled_data = 16'b1011001001001001;
				18'b010010010010011100: oled_data = 16'b1010101000001000;
				18'b010010010100011100: oled_data = 16'b1011101001001001;
				18'b010010010110011100: oled_data = 16'b1011001001001001;
				18'b010010011000011100: oled_data = 16'b1010000111101000;
				18'b010010011010011100: oled_data = 16'b1010000111000111;
				18'b010010011100011100: oled_data = 16'b1011001001001001;
				18'b010010011110011100: oled_data = 16'b1011001000101000;
				18'b010010100000011100: oled_data = 16'b1011001000101001;
				18'b010010100010011100: oled_data = 16'b1011001000101000;
				18'b010010100100011100: oled_data = 16'b1011001000101000;
				18'b010010100110011100: oled_data = 16'b1010101000101000;
				18'b010000011000011101: oled_data = 16'b0101101011001001;
				18'b010000011010011101: oled_data = 16'b1001010001001100;
				18'b010000011100011101: oled_data = 16'b1011010100110000;
				18'b010000011110011101: oled_data = 16'b1010110111110001;
				18'b010000100000011101: oled_data = 16'b1010010111110011;
				18'b010000100010011101: oled_data = 16'b1001010111110100;
				18'b010000100100011101: oled_data = 16'b1001011000010100;
				18'b010000100110011101: oled_data = 16'b1000110110010011;
				18'b010000101000011101: oled_data = 16'b1011110000010011;
				18'b010000101010011101: oled_data = 16'b1101110011010101;
				18'b010000101100011101: oled_data = 16'b1101110011010110;
				18'b010000101110011101: oled_data = 16'b1110010011110110;
				18'b010000110000011101: oled_data = 16'b1101010001110100;
				18'b010000110010011101: oled_data = 16'b1101110010110101;
				18'b010000110100011101: oled_data = 16'b1101110011010110;
				18'b010000110110011101: oled_data = 16'b1101010001110100;
				18'b010000111000011101: oled_data = 16'b1101110011010110;
				18'b010000111010011101: oled_data = 16'b1101010001110100;
				18'b010000111100011101: oled_data = 16'b1101010010010101;
				18'b010000111110011101: oled_data = 16'b1101110010110101;
				18'b010001000000011101: oled_data = 16'b1101110011010101;
				18'b010001000010011101: oled_data = 16'b1101110011010101;
				18'b010001000100011101: oled_data = 16'b1101110011010101;
				18'b010001000110011101: oled_data = 16'b1101110011010101;
				18'b010001001000011101: oled_data = 16'b1101010100110110;
				18'b010001001010011101: oled_data = 16'b1110011011111010;
				18'b010001001100011101: oled_data = 16'b1110111100111011;
				18'b010001001110011101: oled_data = 16'b1110011000111001;
				18'b010001010000011101: oled_data = 16'b1101010011010101;
				18'b010001010010011101: oled_data = 16'b1110010010110101;
				18'b010001010100011101: oled_data = 16'b1101110011010101;
				18'b010001010110011101: oled_data = 16'b1100110100010101;
				18'b010001011000011101: oled_data = 16'b1110111011011010;
				18'b010001011010011101: oled_data = 16'b1110011010111010;
				18'b010001011100011101: oled_data = 16'b1101010100010101;
				18'b010001011110011101: oled_data = 16'b1101110010110101;
				18'b010001100000011101: oled_data = 16'b1101110011010101;
				18'b010001100010011101: oled_data = 16'b1101110011010101;
				18'b010001100100011101: oled_data = 16'b1101110011010101;
				18'b010001100110011101: oled_data = 16'b1101110011010101;
				18'b010001101000011101: oled_data = 16'b1101110011010101;
				18'b010001101010011101: oled_data = 16'b1101110011010101;
				18'b010001101100011101: oled_data = 16'b1110010011110110;
				18'b010001101110011101: oled_data = 16'b1000101010101100;
				18'b010001110000011101: oled_data = 16'b0100000111100111;
				18'b010001110010011101: oled_data = 16'b1101011010011001;
				18'b010001110100011101: oled_data = 16'b1110111100111011;
				18'b010001110110011101: oled_data = 16'b1101011001111001;
				18'b010001111000011101: oled_data = 16'b1011010100010100;
				18'b010001111010011101: oled_data = 16'b0111101101001101;
				18'b010001111100011101: oled_data = 16'b1010110100110011;
				18'b010001111110011101: oled_data = 16'b1101010111110111;
				18'b010010000000011101: oled_data = 16'b1101110011110011;
				18'b010010000010011101: oled_data = 16'b1110010011010011;
				18'b010010000100011101: oled_data = 16'b1011101010001010;
				18'b010010000110011101: oled_data = 16'b1011001000101001;
				18'b010010001000011101: oled_data = 16'b1100001011101011;
				18'b010010001010011101: oled_data = 16'b1100001100101100;
				18'b010010001100011101: oled_data = 16'b1011001000101001;
				18'b010010001110011101: oled_data = 16'b1011101001001001;
				18'b010010010000011101: oled_data = 16'b1011001000101000;
				18'b010010010010011101: oled_data = 16'b1011001001001001;
				18'b010010010100011101: oled_data = 16'b1011101001001001;
				18'b010010010110011101: oled_data = 16'b1010001000001000;
				18'b010010011000011101: oled_data = 16'b1001000101100110;
				18'b010010011010011101: oled_data = 16'b1010101000001000;
				18'b010010011100011101: oled_data = 16'b1011001000101001;
				18'b010010011110011101: oled_data = 16'b1011001000101000;
				18'b010010100000011101: oled_data = 16'b1011001000101001;
				18'b010010100010011101: oled_data = 16'b1011001000101000;
				18'b010010100100011101: oled_data = 16'b1011001000101000;
				18'b010010100110011101: oled_data = 16'b1010101000101000;
				18'b010000011000011110: oled_data = 16'b1100110011110001;
				18'b010000011010011110: oled_data = 16'b1100010100001111;
				18'b010000011100011110: oled_data = 16'b1101110111101110;
				18'b010000011110011110: oled_data = 16'b1110011010010001;
				18'b010000100000011110: oled_data = 16'b1101111010110010;
				18'b010000100010011110: oled_data = 16'b1100111000001101;
				18'b010000100100011110: oled_data = 16'b1100010111001010;
				18'b010000100110011110: oled_data = 16'b1100111000001100;
				18'b010000101000011110: oled_data = 16'b1100010001010000;
				18'b010000101010011110: oled_data = 16'b1101010001110100;
				18'b010000101100011110: oled_data = 16'b1101110011010101;
				18'b010000101110011110: oled_data = 16'b1110010011110110;
				18'b010000110000011110: oled_data = 16'b1100110001010100;
				18'b010000110010011110: oled_data = 16'b1101010001110100;
				18'b010000110100011110: oled_data = 16'b1110010011010110;
				18'b010000110110011110: oled_data = 16'b1101010010010100;
				18'b010000111000011110: oled_data = 16'b1101110011010101;
				18'b010000111010011110: oled_data = 16'b1101010001110100;
				18'b010000111100011110: oled_data = 16'b1101110010110101;
				18'b010000111110011110: oled_data = 16'b1101010010010101;
				18'b010001000000011110: oled_data = 16'b1101110011010110;
				18'b010001000010011110: oled_data = 16'b1101110011010101;
				18'b010001000100011110: oled_data = 16'b1101110011010101;
				18'b010001000110011110: oled_data = 16'b1101110011010110;
				18'b010001001000011110: oled_data = 16'b1101010100010101;
				18'b010001001010011110: oled_data = 16'b1110011011111010;
				18'b010001001100011110: oled_data = 16'b1110111100011010;
				18'b010001001110011110: oled_data = 16'b1110111100011011;
				18'b010001010000011110: oled_data = 16'b1110011000011000;
				18'b010001010010011110: oled_data = 16'b1101010010010100;
				18'b010001010100011110: oled_data = 16'b1101010010010100;
				18'b010001010110011110: oled_data = 16'b1101010010110100;
				18'b010001011000011110: oled_data = 16'b1101111001011000;
				18'b010001011010011110: oled_data = 16'b1110111100111011;
				18'b010001011100011110: oled_data = 16'b1110011010011010;
				18'b010001011110011110: oled_data = 16'b1101010100110101;
				18'b010001100000011110: oled_data = 16'b1101110010110101;
				18'b010001100010011110: oled_data = 16'b1110010011010110;
				18'b010001100100011110: oled_data = 16'b1101110011010101;
				18'b010001100110011110: oled_data = 16'b1101110011010101;
				18'b010001101000011110: oled_data = 16'b1101110011010101;
				18'b010001101010011110: oled_data = 16'b1101110011010110;
				18'b010001101100011110: oled_data = 16'b1101010010010100;
				18'b010001101110011110: oled_data = 16'b0101100110101000;
				18'b010001110000011110: oled_data = 16'b0110101101001101;
				18'b010001110010011110: oled_data = 16'b1010110100110100;
				18'b010001110100011110: oled_data = 16'b0110101100001100;
				18'b010001110110011110: oled_data = 16'b0011100110100110;
				18'b010001111000011110: oled_data = 16'b0100000110100111;
				18'b010001111010011110: oled_data = 16'b1000101111001111;
				18'b010001111100011110: oled_data = 16'b1100111000111000;
				18'b010001111110011110: oled_data = 16'b1100110101110101;
				18'b010010000000011110: oled_data = 16'b1110110100010100;
				18'b010010000010011110: oled_data = 16'b1101001111110000;
				18'b010010000100011110: oled_data = 16'b1011001000101001;
				18'b010010000110011110: oled_data = 16'b1011101001001001;
				18'b010010001000011110: oled_data = 16'b1100001100001100;
				18'b010010001010011110: oled_data = 16'b1011101010001010;
				18'b010010001100011110: oled_data = 16'b1011001001001001;
				18'b010010001110011110: oled_data = 16'b1011001001001001;
				18'b010010010000011110: oled_data = 16'b1010101000101000;
				18'b010010010010011110: oled_data = 16'b1011001001001001;
				18'b010010010100011110: oled_data = 16'b1010101000101000;
				18'b010010010110011110: oled_data = 16'b1000100101100110;
				18'b010010011000011110: oled_data = 16'b1001100110100111;
				18'b010010011010011110: oled_data = 16'b1011101010001010;
				18'b010010011100011110: oled_data = 16'b1011101010101010;
				18'b010010011110011110: oled_data = 16'b1011001000101000;
				18'b010010100000011110: oled_data = 16'b1011001000101001;
				18'b010010100010011110: oled_data = 16'b1011001000101000;
				18'b010010100100011110: oled_data = 16'b1011001000101000;
				18'b010010100110011110: oled_data = 16'b1010101000101000;
				18'b010000011000011111: oled_data = 16'b1100110011010001;
				18'b010000011010011111: oled_data = 16'b1101110111110000;
				18'b010000011100011111: oled_data = 16'b1110111011010101;
				18'b010000011110011111: oled_data = 16'b1101111010010100;
				18'b010000100000011111: oled_data = 16'b1101111010010100;
				18'b010000100010011111: oled_data = 16'b1101011000010000;
				18'b010000100100011111: oled_data = 16'b1010110011101001;
				18'b010000100110011111: oled_data = 16'b1100110111001011;
				18'b010000101000011111: oled_data = 16'b1100110011101111;
				18'b010000101010011111: oled_data = 16'b1101110010110101;
				18'b010000101100011111: oled_data = 16'b1101010001110100;
				18'b010000101110011111: oled_data = 16'b1110010011010110;
				18'b010000110000011111: oled_data = 16'b1101010001110100;
				18'b010000110010011111: oled_data = 16'b1100110000110011;
				18'b010000110100011111: oled_data = 16'b1110010011110110;
				18'b010000110110011111: oled_data = 16'b1101010010010101;
				18'b010000111000011111: oled_data = 16'b1101110010110101;
				18'b010000111010011111: oled_data = 16'b1101010010010101;
				18'b010000111100011111: oled_data = 16'b1101110010110101;
				18'b010000111110011111: oled_data = 16'b1101010001110100;
				18'b010001000000011111: oled_data = 16'b1101110011010101;
				18'b010001000010011111: oled_data = 16'b1101110011010101;
				18'b010001000100011111: oled_data = 16'b1101110011010101;
				18'b010001000110011111: oled_data = 16'b1110010011010110;
				18'b010001001000011111: oled_data = 16'b1101010011110101;
				18'b010001001010011111: oled_data = 16'b1110011011111010;
				18'b010001001100011111: oled_data = 16'b1110111100011011;
				18'b010001001110011111: oled_data = 16'b1110011011111010;
				18'b010001010000011111: oled_data = 16'b1101111010011001;
				18'b010001010010011111: oled_data = 16'b1101010110110111;
				18'b010001010100011111: oled_data = 16'b1100110011110101;
				18'b010001010110011111: oled_data = 16'b1101110011010101;
				18'b010001011000011111: oled_data = 16'b1100110100110101;
				18'b010001011010011111: oled_data = 16'b1110111100011011;
				18'b010001011100011111: oled_data = 16'b1110111100011011;
				18'b010001011110011111: oled_data = 16'b1110011010111010;
				18'b010001100000011111: oled_data = 16'b1101010101010110;
				18'b010001100010011111: oled_data = 16'b1101110010110101;
				18'b010001100100011111: oled_data = 16'b1101110011010101;
				18'b010001100110011111: oled_data = 16'b1101110011010101;
				18'b010001101000011111: oled_data = 16'b1101110011010101;
				18'b010001101010011111: oled_data = 16'b1110010011110110;
				18'b010001101100011111: oled_data = 16'b1010101110110000;
				18'b010001101110011111: oled_data = 16'b0100000110000111;
				18'b010001110000011111: oled_data = 16'b0011000101100101;
				18'b010001110010011111: oled_data = 16'b0011000100100100;
				18'b010001110100011111: oled_data = 16'b0100100111100111;
				18'b010001110110011111: oled_data = 16'b1000110000001111;
				18'b010001111000011111: oled_data = 16'b1101011001011000;
				18'b010001111010011111: oled_data = 16'b1111011101011100;
				18'b010001111100011111: oled_data = 16'b1101011001011000;
				18'b010001111110011111: oled_data = 16'b1101010100010011;
				18'b010010000000011111: oled_data = 16'b1110110100010100;
				18'b010010000010011111: oled_data = 16'b1100001100001101;
				18'b010010000100011111: oled_data = 16'b1011001000101001;
				18'b010010000110011111: oled_data = 16'b1011101001001001;
				18'b010010001000011111: oled_data = 16'b1011101010001010;
				18'b010010001010011111: oled_data = 16'b1011001001001001;
				18'b010010001100011111: oled_data = 16'b1011001001001001;
				18'b010010001110011111: oled_data = 16'b1010101000101000;
				18'b010010010000011111: oled_data = 16'b1011001001001001;
				18'b010010010010011111: oled_data = 16'b1011001000101001;
				18'b010010010100011111: oled_data = 16'b1001000110000111;
				18'b010010010110011111: oled_data = 16'b1001000101100110;
				18'b010010011000011111: oled_data = 16'b1011001001001010;
				18'b010010011010011111: oled_data = 16'b1101001111101111;
				18'b010010011100011111: oled_data = 16'b1011101010001010;
				18'b010010011110011111: oled_data = 16'b1011001000101000;
				18'b010010100000011111: oled_data = 16'b1011001000101001;
				18'b010010100010011111: oled_data = 16'b1011001000101000;
				18'b010010100100011111: oled_data = 16'b1011001000101000;
				18'b010010100110011111: oled_data = 16'b1010101000101000;
				18'b010000011000100000: oled_data = 16'b1101010110001100;
				18'b010000011010100000: oled_data = 16'b1100110111001100;
				18'b010000011100100000: oled_data = 16'b1011110101101100;
				18'b010000011110100000: oled_data = 16'b1011010011101001;
				18'b010000100000100000: oled_data = 16'b1011110100001010;
				18'b010000100010100000: oled_data = 16'b1100110110101101;
				18'b010000100100100000: oled_data = 16'b1010110010101000;
				18'b010000100110100000: oled_data = 16'b1011010100101001;
				18'b010000101000100000: oled_data = 16'b1101010101101110;
				18'b010000101010100000: oled_data = 16'b1101110011010101;
				18'b010000101100100000: oled_data = 16'b1101110010110101;
				18'b010000101110100000: oled_data = 16'b1110010011010110;
				18'b010000110000100000: oled_data = 16'b1100110001010011;
				18'b010000110010100000: oled_data = 16'b1100001111110010;
				18'b010000110100100000: oled_data = 16'b1110010011010110;
				18'b010000110110100000: oled_data = 16'b1101110010110101;
				18'b010000111000100000: oled_data = 16'b1101010010010100;
				18'b010000111010100000: oled_data = 16'b1101110010110101;
				18'b010000111100100000: oled_data = 16'b1101110010110101;
				18'b010000111110100000: oled_data = 16'b1101010010010101;
				18'b010001000000100000: oled_data = 16'b1101110010010101;
				18'b010001000010100000: oled_data = 16'b1101110011010110;
				18'b010001000100100000: oled_data = 16'b1101110011010101;
				18'b010001000110100000: oled_data = 16'b1110010011010110;
				18'b010001001000100000: oled_data = 16'b1101010011110101;
				18'b010001001010100000: oled_data = 16'b1110011011111010;
				18'b010001001100100000: oled_data = 16'b1101111010011001;
				18'b010001001110100000: oled_data = 16'b1101011010011000;
				18'b010001010000100000: oled_data = 16'b1110011011111010;
				18'b010001010010100000: oled_data = 16'b1111011101011100;
				18'b010001010100100000: oled_data = 16'b1110011001111010;
				18'b010001010110100000: oled_data = 16'b1101010011110101;
				18'b010001011000100000: oled_data = 16'b1101010011010100;
				18'b010001011010100000: oled_data = 16'b1101111000011000;
				18'b010001011100100000: oled_data = 16'b1110111100011011;
				18'b010001011110100000: oled_data = 16'b1110111100011010;
				18'b010001100000100000: oled_data = 16'b1110011011011010;
				18'b010001100010100000: oled_data = 16'b1101010110110110;
				18'b010001100100100000: oled_data = 16'b1101010011010100;
				18'b010001100110100000: oled_data = 16'b1101110011010101;
				18'b010001101000100000: oled_data = 16'b1110010011010110;
				18'b010001101010100000: oled_data = 16'b1101110011010110;
				18'b010001101100100000: oled_data = 16'b1000101010101100;
				18'b010001101110100000: oled_data = 16'b0101001000101001;
				18'b010001110000100000: oled_data = 16'b0111101110101110;
				18'b010001110010100000: oled_data = 16'b1011110101110101;
				18'b010001110100100000: oled_data = 16'b1101111010111010;
				18'b010001110110100000: oled_data = 16'b1110111100111011;
				18'b010001111000100000: oled_data = 16'b1110111100111011;
				18'b010001111010100000: oled_data = 16'b1110011011111010;
				18'b010001111100100000: oled_data = 16'b1101111000111000;
				18'b010001111110100000: oled_data = 16'b1101110011110100;
				18'b010010000000100000: oled_data = 16'b1110010011010011;
				18'b010010000010100000: oled_data = 16'b1011001001101010;
				18'b010010000100100000: oled_data = 16'b1011001000101001;
				18'b010010000110100000: oled_data = 16'b1011001001001001;
				18'b010010001000100000: oled_data = 16'b1011001001001001;
				18'b010010001010100000: oled_data = 16'b1011001001001001;
				18'b010010001100100000: oled_data = 16'b1011001001001001;
				18'b010010001110100000: oled_data = 16'b1010101000101001;
				18'b010010010000100000: oled_data = 16'b1011001001001001;
				18'b010010010010100000: oled_data = 16'b1001100110100111;
				18'b010010010100100000: oled_data = 16'b1000100101000110;
				18'b010010010110100000: oled_data = 16'b1010000111001000;
				18'b010010011000100000: oled_data = 16'b1100101101001101;
				18'b010010011010100000: oled_data = 16'b1100001100001100;
				18'b010010011100100000: oled_data = 16'b1011001000101000;
				18'b010010011110100000: oled_data = 16'b1011001000101001;
				18'b010010100000100000: oled_data = 16'b1011001000101001;
				18'b010010100010100000: oled_data = 16'b1011001000101000;
				18'b010010100100100000: oled_data = 16'b1011001000101000;
				18'b010010100110100000: oled_data = 16'b1010101000101000;
				18'b010000011000100001: oled_data = 16'b1101010111101011;
				18'b010000011010100001: oled_data = 16'b1011010011100111;
				18'b010000011100100001: oled_data = 16'b1010110010100111;
				18'b010000011110100001: oled_data = 16'b1010110010100111;
				18'b010000100000100001: oled_data = 16'b1010110011001000;
				18'b010000100010100001: oled_data = 16'b1100010101101011;
				18'b010000100100100001: oled_data = 16'b1010110011001000;
				18'b010000100110100001: oled_data = 16'b1010110011001000;
				18'b010000101000100001: oled_data = 16'b1101010110001101;
				18'b010000101010100001: oled_data = 16'b1101110011010101;
				18'b010000101100100001: oled_data = 16'b1101010010010100;
				18'b010000101110100001: oled_data = 16'b1101110011010101;
				18'b010000110000100001: oled_data = 16'b1100110000110011;
				18'b010000110010100001: oled_data = 16'b1011101110110001;
				18'b010000110100100001: oled_data = 16'b1101110011010110;
				18'b010000110110100001: oled_data = 16'b1101110011010101;
				18'b010000111000100001: oled_data = 16'b1101010001110100;
				18'b010000111010100001: oled_data = 16'b1101110010110101;
				18'b010000111100100001: oled_data = 16'b1101010001110100;
				18'b010000111110100001: oled_data = 16'b1101110011010101;
				18'b010001000000100001: oled_data = 16'b1101010010010100;
				18'b010001000010100001: oled_data = 16'b1101110011010101;
				18'b010001000100100001: oled_data = 16'b1101110011010101;
				18'b010001000110100001: oled_data = 16'b1110010011010110;
				18'b010001001000100001: oled_data = 16'b1101010011110101;
				18'b010001001010100001: oled_data = 16'b1101011001011000;
				18'b010001001100100001: oled_data = 16'b1101111010111001;
				18'b010001001110100001: oled_data = 16'b1110011100011011;
				18'b010001010000100001: oled_data = 16'b1110111100011011;
				18'b010001010010100001: oled_data = 16'b1110111100011011;
				18'b010001010100100001: oled_data = 16'b1111011100111100;
				18'b010001010110100001: oled_data = 16'b1110111010011010;
				18'b010001011000100001: oled_data = 16'b1101010101010110;
				18'b010001011010100001: oled_data = 16'b1100010011110100;
				18'b010001011100100001: oled_data = 16'b1110011010111010;
				18'b010001011110100001: oled_data = 16'b1110111100011010;
				18'b010001100000100001: oled_data = 16'b1110111100011010;
				18'b010001100010100001: oled_data = 16'b1110111100011010;
				18'b010001100100100001: oled_data = 16'b1101111000010111;
				18'b010001100110100001: oled_data = 16'b1100110011110101;
				18'b010001101000100001: oled_data = 16'b1101010010110101;
				18'b010001101010100001: oled_data = 16'b1101110011010101;
				18'b010001101100100001: oled_data = 16'b1100010000110011;
				18'b010001101110100001: oled_data = 16'b1100110110110110;
				18'b010001110000100001: oled_data = 16'b1111011101111100;
				18'b010001110010100001: oled_data = 16'b1111011100111011;
				18'b010001110100100001: oled_data = 16'b1110111100011011;
				18'b010001110110100001: oled_data = 16'b1110011100011010;
				18'b010001111000100001: oled_data = 16'b1110011100011010;
				18'b010001111010100001: oled_data = 16'b1101111010011001;
				18'b010001111100100001: oled_data = 16'b1101111000010111;
				18'b010001111110100001: oled_data = 16'b1110010100010100;
				18'b010010000000100001: oled_data = 16'b1101110001110001;
				18'b010010000010100001: oled_data = 16'b1011001000101001;
				18'b010010000100100001: oled_data = 16'b1011001001001001;
				18'b010010000110100001: oled_data = 16'b1011001001001001;
				18'b010010001000100001: oled_data = 16'b1011001001001001;
				18'b010010001010100001: oled_data = 16'b1011001001001001;
				18'b010010001100100001: oled_data = 16'b1010101000101001;
				18'b010010001110100001: oled_data = 16'b1011001001001001;
				18'b010010010000100001: oled_data = 16'b1010000111101000;
				18'b010010010010100001: oled_data = 16'b1000100101000110;
				18'b010010010100100001: oled_data = 16'b1001100110000111;
				18'b010010010110100001: oled_data = 16'b1011001000101001;
				18'b010010011000100001: oled_data = 16'b1011101010001010;
				18'b010010011010100001: oled_data = 16'b1011001001001001;
				18'b010010011100100001: oled_data = 16'b1011001000101001;
				18'b010010011110100001: oled_data = 16'b1011001000101001;
				18'b010010100000100001: oled_data = 16'b1011001000101001;
				18'b010010100010100001: oled_data = 16'b1011001000101000;
				18'b010010100100100001: oled_data = 16'b1011001000101000;
				18'b010010100110100001: oled_data = 16'b1010101000101000;
				18'b010000011000100010: oled_data = 16'b1100010110001011;
				18'b010000011010100010: oled_data = 16'b1011010011101000;
				18'b010000011100100010: oled_data = 16'b1010110010100111;
				18'b010000011110100010: oled_data = 16'b1010110010100111;
				18'b010000100000100010: oled_data = 16'b1010110010100111;
				18'b010000100010100010: oled_data = 16'b1011110100101010;
				18'b010000100100100010: oled_data = 16'b1010110011001001;
				18'b010000100110100010: oled_data = 16'b1010110011001000;
				18'b010000101000100010: oled_data = 16'b1100110110101100;
				18'b010000101010100010: oled_data = 16'b1101110011010101;
				18'b010000101100100010: oled_data = 16'b1100110000110011;
				18'b010000101110100010: oled_data = 16'b1011101111010001;
				18'b010000110000100010: oled_data = 16'b1011101111010001;
				18'b010000110010100010: oled_data = 16'b1011101110110001;
				18'b010000110100100010: oled_data = 16'b1101110011010101;
				18'b010000110110100010: oled_data = 16'b1101110011010110;
				18'b010000111000100010: oled_data = 16'b1101010010010100;
				18'b010000111010100010: oled_data = 16'b1101010010010100;
				18'b010000111100100010: oled_data = 16'b1101010001110100;
				18'b010000111110100010: oled_data = 16'b1101110011010110;
				18'b010001000000100010: oled_data = 16'b1101010001110100;
				18'b010001000010100010: oled_data = 16'b1101110010110101;
				18'b010001000100100010: oled_data = 16'b1101110011010110;
				18'b010001000110100010: oled_data = 16'b1101110011010110;
				18'b010001001000100010: oled_data = 16'b1101110100010110;
				18'b010001001010100010: oled_data = 16'b1110011011111011;
				18'b010001001100100010: oled_data = 16'b1110111100011011;
				18'b010001001110100010: oled_data = 16'b1110111100011011;
				18'b010001010000100010: oled_data = 16'b1110111100011011;
				18'b010001010010100010: oled_data = 16'b1110111100011010;
				18'b010001010100100010: oled_data = 16'b1110111100011010;
				18'b010001010110100010: oled_data = 16'b1110111100011011;
				18'b010001011000100010: oled_data = 16'b1110111011111010;
				18'b010001011010100010: oled_data = 16'b1101010111010111;
				18'b010001011100100010: oled_data = 16'b1100110110110110;
				18'b010001011110100010: oled_data = 16'b1110111100011010;
				18'b010001100000100010: oled_data = 16'b1110011100011010;
				18'b010001100010100010: oled_data = 16'b1110011100011010;
				18'b010001100100100010: oled_data = 16'b1110011100111010;
				18'b010001100110100010: oled_data = 16'b1110011010111010;
				18'b010001101000100010: oled_data = 16'b1100110110010110;
				18'b010001101010100010: oled_data = 16'b1101010011110101;
				18'b010001101100100010: oled_data = 16'b1101010010110101;
				18'b010001101110100010: oled_data = 16'b1101111001011000;
				18'b010001110000100010: oled_data = 16'b1110111100011010;
				18'b010001110010100010: oled_data = 16'b1110111100011010;
				18'b010001110100100010: oled_data = 16'b1110111100011010;
				18'b010001110110100010: oled_data = 16'b1110111100011010;
				18'b010001111000100010: oled_data = 16'b1101111011011001;
				18'b010001111010100010: oled_data = 16'b1110011011011010;
				18'b010001111100100010: oled_data = 16'b1101110110110110;
				18'b010001111110100010: oled_data = 16'b1110010100010100;
				18'b010010000000100010: oled_data = 16'b1100101111001111;
				18'b010010000010100010: oled_data = 16'b1011001000001000;
				18'b010010000100100010: oled_data = 16'b1011101001001001;
				18'b010010000110100010: oled_data = 16'b1011001001001001;
				18'b010010001000100010: oled_data = 16'b1011001001001001;
				18'b010010001010100010: oled_data = 16'b1011001001001001;
				18'b010010001100100010: oled_data = 16'b1010101000101000;
				18'b010010001110100010: oled_data = 16'b1011001001001001;
				18'b010010010000100010: oled_data = 16'b1001000101100111;
				18'b010010010010100010: oled_data = 16'b1000100101000110;
				18'b010010010100100010: oled_data = 16'b1010101000001000;
				18'b010010010110100010: oled_data = 16'b1011001001001001;
				18'b010010011000100010: oled_data = 16'b1011001001001001;
				18'b010010011010100010: oled_data = 16'b1011001001001001;
				18'b010010011100100010: oled_data = 16'b1011001001001001;
				18'b010010011110100010: oled_data = 16'b1011001001001001;
				18'b010010100000100010: oled_data = 16'b1011001000101001;
				18'b010010100010100010: oled_data = 16'b1011001000101000;
				18'b010010100100100010: oled_data = 16'b1010101000101000;
				18'b010010100110100010: oled_data = 16'b1010101000101000;
				18'b010000011000100011: oled_data = 16'b1011010100101011;
				18'b010000011010100011: oled_data = 16'b1011010100001000;
				18'b010000011100100011: oled_data = 16'b1010110010100111;
				18'b010000011110100011: oled_data = 16'b1010110010100111;
				18'b010000100000100011: oled_data = 16'b1010110010100111;
				18'b010000100010100011: oled_data = 16'b1011010011101000;
				18'b010000100100100011: oled_data = 16'b1010110011001000;
				18'b010000100110100011: oled_data = 16'b1010110011000111;
				18'b010000101000100011: oled_data = 16'b1101010111001100;
				18'b010000101010100011: oled_data = 16'b1101110011110101;
				18'b010000101100100011: oled_data = 16'b1101110010110101;
				18'b010000101110100011: oled_data = 16'b1011101111010001;
				18'b010000110000100011: oled_data = 16'b1011001110010000;
				18'b010000110010100011: oled_data = 16'b1011001101110000;
				18'b010000110100100011: oled_data = 16'b1101110010110101;
				18'b010000110110100011: oled_data = 16'b1101110011010110;
				18'b010000111000100011: oled_data = 16'b1101110010110101;
				18'b010000111010100011: oled_data = 16'b1101010001110100;
				18'b010000111100100011: oled_data = 16'b1101010001110100;
				18'b010000111110100011: oled_data = 16'b1101110011010101;
				18'b010001000000100011: oled_data = 16'b1101110010110101;
				18'b010001000010100011: oled_data = 16'b1101010010010100;
				18'b010001000100100011: oled_data = 16'b1101110011010101;
				18'b010001000110100011: oled_data = 16'b1101110011010101;
				18'b010001001000100011: oled_data = 16'b1101010101010110;
				18'b010001001010100011: oled_data = 16'b1110111100011011;
				18'b010001001100100011: oled_data = 16'b1110111100011011;
				18'b010001001110100011: oled_data = 16'b1110111100111011;
				18'b010001010000100011: oled_data = 16'b1110111100111011;
				18'b010001010010100011: oled_data = 16'b1111011100111011;
				18'b010001010100100011: oled_data = 16'b1111011101011011;
				18'b010001010110100011: oled_data = 16'b1111011100111100;
				18'b010001011000100011: oled_data = 16'b1111011100111011;
				18'b010001011010100011: oled_data = 16'b1111011100011011;
				18'b010001011100100011: oled_data = 16'b1101111001011000;
				18'b010001011110100011: oled_data = 16'b1101111010011001;
				18'b010001100000100011: oled_data = 16'b1101111010111001;
				18'b010001100010100011: oled_data = 16'b1110011100011010;
				18'b010001100100100011: oled_data = 16'b1110011100011010;
				18'b010001100110100011: oled_data = 16'b1110011100011011;
				18'b010001101000100011: oled_data = 16'b1110011011111010;
				18'b010001101010100011: oled_data = 16'b1110011001111010;
				18'b010001101100100011: oled_data = 16'b1101010110010111;
				18'b010001101110100011: oled_data = 16'b1110011010011001;
				18'b010001110000100011: oled_data = 16'b1110111100011010;
				18'b010001110010100011: oled_data = 16'b1110111100011010;
				18'b010001110100100011: oled_data = 16'b1110111100011010;
				18'b010001110110100011: oled_data = 16'b1110011011111010;
				18'b010001111000100011: oled_data = 16'b1101111010011001;
				18'b010001111010100011: oled_data = 16'b1110111100011011;
				18'b010001111100100011: oled_data = 16'b1101110110010110;
				18'b010001111110100011: oled_data = 16'b1110010100010100;
				18'b010010000000100011: oled_data = 16'b1100001100101100;
				18'b010010000010100011: oled_data = 16'b1011001000101000;
				18'b010010000100100011: oled_data = 16'b1011101001001001;
				18'b010010000110100011: oled_data = 16'b1011001001001001;
				18'b010010001000100011: oled_data = 16'b1011001001001001;
				18'b010010001010100011: oled_data = 16'b1011001000101001;
				18'b010010001100100011: oled_data = 16'b1010101000101001;
				18'b010010001110100011: oled_data = 16'b1010000111101000;
				18'b010010010000100011: oled_data = 16'b1000100101000110;
				18'b010010010010100011: oled_data = 16'b1001100111001000;
				18'b010010010100100011: oled_data = 16'b1011001001001001;
				18'b010010010110100011: oled_data = 16'b1011001001001001;
				18'b010010011000100011: oled_data = 16'b1011001001001001;
				18'b010010011010100011: oled_data = 16'b1011001001001001;
				18'b010010011100100011: oled_data = 16'b1011001000101001;
				18'b010010011110100011: oled_data = 16'b1011001000101001;
				18'b010010100000100011: oled_data = 16'b1011001000101001;
				18'b010010100010100011: oled_data = 16'b1011001000101000;
				18'b010010100100100011: oled_data = 16'b1010101000101000;
				18'b010010100110100011: oled_data = 16'b1010101000101000;
				18'b010000011000100100: oled_data = 16'b1010010011001010;
				18'b010000011010100100: oled_data = 16'b1100010101101001;
				18'b010000011100100100: oled_data = 16'b1010110010100111;
				18'b010000011110100100: oled_data = 16'b1010110010100111;
				18'b010000100000100100: oled_data = 16'b1010110010100111;
				18'b010000100010100100: oled_data = 16'b1010110010100111;
				18'b010000100100100100: oled_data = 16'b1010110010100111;
				18'b010000100110100100: oled_data = 16'b1011010011101000;
				18'b010000101000100100: oled_data = 16'b1101010111101101;
				18'b010000101010100100: oled_data = 16'b1101110011110100;
				18'b010000101100100100: oled_data = 16'b1110010011010110;
				18'b010000101110100100: oled_data = 16'b1101010010010100;
				18'b010000110000100100: oled_data = 16'b1011001111010001;
				18'b010000110010100100: oled_data = 16'b1010101101110000;
				18'b010000110100100100: oled_data = 16'b1101010010010100;
				18'b010000110110100100: oled_data = 16'b1101110011010110;
				18'b010000111000100100: oled_data = 16'b1101110011010110;
				18'b010000111010100100: oled_data = 16'b1101110010010101;
				18'b010000111100100100: oled_data = 16'b1101010001110100;
				18'b010000111110100100: oled_data = 16'b1101110011010101;
				18'b010001000000100100: oled_data = 16'b1101110011010101;
				18'b010001000010100100: oled_data = 16'b1101110010110101;
				18'b010001000100100100: oled_data = 16'b1101010010010100;
				18'b010001000110100100: oled_data = 16'b1110010011110101;
				18'b010001001000100100: oled_data = 16'b1101110110110110;
				18'b010001001010100100: oled_data = 16'b1110111011111011;
				18'b010001001100100100: oled_data = 16'b1101111010111010;
				18'b010001001110100100: oled_data = 16'b1101011001111001;
				18'b010001010000100100: oled_data = 16'b1100110111110111;
				18'b010001010010100100: oled_data = 16'b1011010101010100;
				18'b010001010100100100: oled_data = 16'b1001110010110010;
				18'b010001010110100100: oled_data = 16'b1000110000110000;
				18'b010001011000100100: oled_data = 16'b0111001101101100;
				18'b010001011010100100: oled_data = 16'b0110001011001011;
				18'b010001011100100100: oled_data = 16'b0101101001101001;
				18'b010001011110100100: oled_data = 16'b0100100111100111;
				18'b010001100000100100: oled_data = 16'b1001010001110000;
				18'b010001100010100100: oled_data = 16'b1110111100111011;
				18'b010001100100100100: oled_data = 16'b1110011100011010;
				18'b010001100110100100: oled_data = 16'b1110011100011010;
				18'b010001101000100100: oled_data = 16'b1110011100011010;
				18'b010001101010100100: oled_data = 16'b1110011100011010;
				18'b010001101100100100: oled_data = 16'b1110111100011010;
				18'b010001101110100100: oled_data = 16'b1110111100011010;
				18'b010001110000100100: oled_data = 16'b1110111011111010;
				18'b010001110010100100: oled_data = 16'b1110111100011010;
				18'b010001110100100100: oled_data = 16'b1110111100011011;
				18'b010001110110100100: oled_data = 16'b1101111010111010;
				18'b010001111000100100: oled_data = 16'b1110111100011011;
				18'b010001111010100100: oled_data = 16'b1110111011111010;
				18'b010001111100100100: oled_data = 16'b1101010101010101;
				18'b010001111110100100: oled_data = 16'b1110110011110011;
				18'b010010000000100100: oled_data = 16'b1011001010101011;
				18'b010010000010100100: oled_data = 16'b1011001000101001;
				18'b010010000100100100: oled_data = 16'b1011001001001001;
				18'b010010000110100100: oled_data = 16'b1011001001001001;
				18'b010010001000100100: oled_data = 16'b1011001001001001;
				18'b010010001010100100: oled_data = 16'b1010101000101000;
				18'b010010001100100100: oled_data = 16'b1011001000101001;
				18'b010010001110100100: oled_data = 16'b1001000101100110;
				18'b010010010000100100: oled_data = 16'b1001000101100111;
				18'b010010010010100100: oled_data = 16'b1011001000101001;
				18'b010010010100100100: oled_data = 16'b1011001001001001;
				18'b010010010110100100: oled_data = 16'b1011001000101001;
				18'b010010011000100100: oled_data = 16'b1011001001001001;
				18'b010010011010100100: oled_data = 16'b1011001001001001;
				18'b010010011100100100: oled_data = 16'b1011001001001001;
				18'b010010011110100100: oled_data = 16'b1011001001001001;
				18'b010010100000100100: oled_data = 16'b1011001000101001;
				18'b010010100010100100: oled_data = 16'b1011001000101000;
				18'b010010100100100100: oled_data = 16'b1010101000101000;
				18'b010010100110100100: oled_data = 16'b1010101000101000;
				18'b010000011000100101: oled_data = 16'b1000001111001001;
				18'b010000011010100101: oled_data = 16'b1101011000001011;
				18'b010000011100100101: oled_data = 16'b1011010100001000;
				18'b010000011110100101: oled_data = 16'b1010110010100111;
				18'b010000100000100101: oled_data = 16'b1010110010100111;
				18'b010000100010100101: oled_data = 16'b1010110010100111;
				18'b010000100100100101: oled_data = 16'b1010110011000111;
				18'b010000100110100101: oled_data = 16'b1100110110101010;
				18'b010000101000100101: oled_data = 16'b1101110111101101;
				18'b010000101010100101: oled_data = 16'b1101110011110101;
				18'b010000101100100101: oled_data = 16'b1101110011010101;
				18'b010000101110100101: oled_data = 16'b1101010101010110;
				18'b010000110000100101: oled_data = 16'b1101111001011001;
				18'b010000110010100101: oled_data = 16'b1100110101010101;
				18'b010000110100100101: oled_data = 16'b1101010010010100;
				18'b010000110110100101: oled_data = 16'b1101110011010101;
				18'b010000111000100101: oled_data = 16'b1101110011010101;
				18'b010000111010100101: oled_data = 16'b1101110011010101;
				18'b010000111100100101: oled_data = 16'b1100110001010011;
				18'b010000111110100101: oled_data = 16'b1101110010110101;
				18'b010001000000100101: oled_data = 16'b1101110011010110;
				18'b010001000010100101: oled_data = 16'b1110010011010110;
				18'b010001000100100101: oled_data = 16'b1100010000010010;
				18'b010001000110100101: oled_data = 16'b1000101010001100;
				18'b010001001000100101: oled_data = 16'b0110101010001010;
				18'b010001001010100101: oled_data = 16'b0101101001101001;
				18'b010001001100100101: oled_data = 16'b0100101000000111;
				18'b010001001110100101: oled_data = 16'b0011100110100110;
				18'b010001010000100101: oled_data = 16'b0011000101100101;
				18'b010001010010100101: oled_data = 16'b0010100100000100;
				18'b010001010100100101: oled_data = 16'b0010100100000100;
				18'b010001010110100101: oled_data = 16'b0010100100100100;
				18'b010001011000100101: oled_data = 16'b0011100110100110;
				18'b010001011010100101: oled_data = 16'b0011000101100101;
				18'b010001011100100101: oled_data = 16'b0011000100100100;
				18'b010001011110100101: oled_data = 16'b0101101001101001;
				18'b010001100000100101: oled_data = 16'b1101011001111000;
				18'b010001100010100101: oled_data = 16'b1110111100011010;
				18'b010001100100100101: oled_data = 16'b1110011100011010;
				18'b010001100110100101: oled_data = 16'b1110011100011010;
				18'b010001101000100101: oled_data = 16'b1110011100011010;
				18'b010001101010100101: oled_data = 16'b1110011100011010;
				18'b010001101100100101: oled_data = 16'b1110011100011010;
				18'b010001101110100101: oled_data = 16'b1110111011111011;
				18'b010001110000100101: oled_data = 16'b1110111011111010;
				18'b010001110010100101: oled_data = 16'b1110111100011010;
				18'b010001110100100101: oled_data = 16'b1101111010111001;
				18'b010001110110100101: oled_data = 16'b1110011011011010;
				18'b010001111000100101: oled_data = 16'b1110111100011011;
				18'b010001111010100101: oled_data = 16'b1110011010111010;
				18'b010001111100100101: oled_data = 16'b1101110100010100;
				18'b010001111110100101: oled_data = 16'b1110010011010011;
				18'b010010000000100101: oled_data = 16'b1011001001101001;
				18'b010010000010100101: oled_data = 16'b1011001001001001;
				18'b010010000100100101: oled_data = 16'b1011001001001001;
				18'b010010000110100101: oled_data = 16'b1011001001001001;
				18'b010010001000100101: oled_data = 16'b1011101010101010;
				18'b010010001010100101: oled_data = 16'b1011001010001001;
				18'b010010001100100101: oled_data = 16'b1010000111100111;
				18'b010010001110100101: oled_data = 16'b1000100101000110;
				18'b010010010000100101: oled_data = 16'b1010000111101001;
				18'b010010010010100101: oled_data = 16'b1011001001001001;
				18'b010010010100100101: oled_data = 16'b1011001000101000;
				18'b010010010110100101: oled_data = 16'b1011101110101111;
				18'b010010011000100101: oled_data = 16'b1011001010101011;
				18'b010010011010100101: oled_data = 16'b1011001001001001;
				18'b010010011100100101: oled_data = 16'b1011101010001010;
				18'b010010011110100101: oled_data = 16'b1011001001001001;
				18'b010010100000100101: oled_data = 16'b1011001000101001;
				18'b010010100010100101: oled_data = 16'b1011001000101000;
				18'b010010100100100101: oled_data = 16'b1010101000101000;
				18'b010010100110100101: oled_data = 16'b1010101000101000;
				18'b010000011000100110: oled_data = 16'b0101001010000110;
				18'b010000011010100110: oled_data = 16'b1100111000001011;
				18'b010000011100100110: oled_data = 16'b1101011001001011;
				18'b010000011110100110: oled_data = 16'b1100010111001001;
				18'b010000100000100110: oled_data = 16'b1100110110101001;
				18'b010000100010100110: oled_data = 16'b1100010110001001;
				18'b010000100100100110: oled_data = 16'b1100110111101011;
				18'b010000100110100110: oled_data = 16'b1101010110101100;
				18'b010000101000100110: oled_data = 16'b1101010100010000;
				18'b010000101010100110: oled_data = 16'b1101110011010101;
				18'b010000101100100110: oled_data = 16'b1101110011010101;
				18'b010000101110100110: oled_data = 16'b1101111000111000;
				18'b010000110000100110: oled_data = 16'b1101011001011000;
				18'b010000110010100110: oled_data = 16'b1101110111111000;
				18'b010000110100100110: oled_data = 16'b1101010011010100;
				18'b010000110110100110: oled_data = 16'b1101110010110101;
				18'b010000111000100110: oled_data = 16'b1101110011010101;
				18'b010000111010100110: oled_data = 16'b1101110011010110;
				18'b010000111100100110: oled_data = 16'b1101010010010100;
				18'b010000111110100110: oled_data = 16'b1101010001110100;
				18'b010001000000100110: oled_data = 16'b1101110011010110;
				18'b010001000010100110: oled_data = 16'b1101110011010101;
				18'b010001000100100110: oled_data = 16'b1101110011010101;
				18'b010001000110100110: oled_data = 16'b1000001100001101;
				18'b010001001000100110: oled_data = 16'b0100101000101000;
				18'b010001001010100110: oled_data = 16'b0101001001001000;
				18'b010001001100100110: oled_data = 16'b0110001011001010;
				18'b010001001110100110: oled_data = 16'b0110001100101100;
				18'b010001010000100110: oled_data = 16'b0110101100101100;
				18'b010001010010100110: oled_data = 16'b1000001111101110;
				18'b010001010100100110: oled_data = 16'b1001110010110010;
				18'b010001010110100110: oled_data = 16'b1011110110010110;
				18'b010001011000100110: oled_data = 16'b0111001101001100;
				18'b010001011010100110: oled_data = 16'b0010100101000100;
				18'b010001011100100110: oled_data = 16'b0100101000000111;
				18'b010001011110100110: oled_data = 16'b1100111000111000;
				18'b010001100000100110: oled_data = 16'b1110111100111011;
				18'b010001100010100110: oled_data = 16'b1110111100011010;
				18'b010001100100100110: oled_data = 16'b1110111100011010;
				18'b010001100110100110: oled_data = 16'b1110111100011010;
				18'b010001101000100110: oled_data = 16'b1110111100011010;
				18'b010001101010100110: oled_data = 16'b1110111100011011;
				18'b010001101100100110: oled_data = 16'b1110111100011010;
				18'b010001101110100110: oled_data = 16'b1110111100011011;
				18'b010001110000100110: oled_data = 16'b1110111100011011;
				18'b010001110010100110: oled_data = 16'b1110011011111010;
				18'b010001110100100110: oled_data = 16'b1101111010011001;
				18'b010001110110100110: oled_data = 16'b1110111100011010;
				18'b010001111000100110: oled_data = 16'b1110111100011011;
				18'b010001111010100110: oled_data = 16'b1110011010011001;
				18'b010001111100100110: oled_data = 16'b1101110011110100;
				18'b010001111110100110: oled_data = 16'b1101110001110001;
				18'b010010000000100110: oled_data = 16'b1010101000101001;
				18'b010010000010100110: oled_data = 16'b1011001001001001;
				18'b010010000100100110: oled_data = 16'b1011001010101010;
				18'b010010000110100110: oled_data = 16'b1101010000110000;
				18'b010010001000100110: oled_data = 16'b1110010010110011;
				18'b010010001010100110: oled_data = 16'b1100101110101111;
				18'b010010001100100110: oled_data = 16'b1010000111101000;
				18'b010010001110100110: oled_data = 16'b1001100110000111;
				18'b010010010000100110: oled_data = 16'b1011001001101010;
				18'b010010010010100110: oled_data = 16'b1011001001001001;
				18'b010010010100100110: oled_data = 16'b1011001001101010;
				18'b010010010110100110: oled_data = 16'b1100011000111001;
				18'b010010011000100110: oled_data = 16'b1011001111110000;
				18'b010010011010100110: oled_data = 16'b1011001000001000;
				18'b010010011100100110: oled_data = 16'b1011001001001001;
				18'b010010011110100110: oled_data = 16'b1011001000101001;
				18'b010010100000100110: oled_data = 16'b1011001000101001;
				18'b010010100010100110: oled_data = 16'b1011001000101000;
				18'b010010100100100110: oled_data = 16'b1010101000101000;
				18'b010010100110100110: oled_data = 16'b1010101000101000;
				18'b010000011000100111: oled_data = 16'b0010000100100100;
				18'b010000011010100111: oled_data = 16'b0110001010100110;
				18'b010000011100100111: oled_data = 16'b1000110000101000;
				18'b010000011110100111: oled_data = 16'b1010010011101011;
				18'b010000100000100111: oled_data = 16'b1011010100101101;
				18'b010000100010100111: oled_data = 16'b1011110011101110;
				18'b010000100100100111: oled_data = 16'b1100010001101111;
				18'b010000100110100111: oled_data = 16'b1011001110010000;
				18'b010000101000100111: oled_data = 16'b1100110001010100;
				18'b010000101010100111: oled_data = 16'b1110010011010110;
				18'b010000101100100111: oled_data = 16'b1101110010110101;
				18'b010000101110100111: oled_data = 16'b1110011001111001;
				18'b010000110000100111: oled_data = 16'b1110011011011010;
				18'b010000110010100111: oled_data = 16'b1101010111110111;
				18'b010000110100100111: oled_data = 16'b1100110010110100;
				18'b010000110110100111: oled_data = 16'b1101110011010101;
				18'b010000111000100111: oled_data = 16'b1101110011010101;
				18'b010000111010100111: oled_data = 16'b1101110011010101;
				18'b010000111100100111: oled_data = 16'b1101110011010101;
				18'b010000111110100111: oled_data = 16'b1101110010110101;
				18'b010001000000100111: oled_data = 16'b1101110011010101;
				18'b010001000010100111: oled_data = 16'b1101110011010101;
				18'b010001000100100111: oled_data = 16'b1101110011010101;
				18'b010001000110100111: oled_data = 16'b1100110101010110;
				18'b010001001000100111: oled_data = 16'b1110011011011010;
				18'b010001001010100111: oled_data = 16'b1110011011111010;
				18'b010001001100100111: oled_data = 16'b1110011100011011;
				18'b010001001110100111: oled_data = 16'b1110011100111011;
				18'b010001010000100111: oled_data = 16'b1110011100111011;
				18'b010001010010100111: oled_data = 16'b1110111100111011;
				18'b010001010100100111: oled_data = 16'b1111011101011100;
				18'b010001010110100111: oled_data = 16'b1010010011010011;
				18'b010001011000100111: oled_data = 16'b0011100101100101;
				18'b010001011010100111: oled_data = 16'b0011100110100110;
				18'b010001011100100111: oled_data = 16'b1011110110010101;
				18'b010001011110100111: oled_data = 16'b1110111100111100;
				18'b010001100000100111: oled_data = 16'b1110111100011011;
				18'b010001100010100111: oled_data = 16'b1110111100011010;
				18'b010001100100100111: oled_data = 16'b1110111100011010;
				18'b010001100110100111: oled_data = 16'b1110111100011010;
				18'b010001101000100111: oled_data = 16'b1110111100011010;
				18'b010001101010100111: oled_data = 16'b1110111100011011;
				18'b010001101100100111: oled_data = 16'b1110111100011010;
				18'b010001101110100111: oled_data = 16'b1110111100011011;
				18'b010001110000100111: oled_data = 16'b1110011100011010;
				18'b010001110010100111: oled_data = 16'b1101111010011001;
				18'b010001110100100111: oled_data = 16'b1110011011111010;
				18'b010001110110100111: oled_data = 16'b1110111100011010;
				18'b010001111000100111: oled_data = 16'b1110011011011010;
				18'b010001111010100111: oled_data = 16'b1100110100110101;
				18'b010001111100100111: oled_data = 16'b1101110011110100;
				18'b010001111110100111: oled_data = 16'b1101010000010000;
				18'b010010000000100111: oled_data = 16'b1010101000101000;
				18'b010010000010100111: oled_data = 16'b1011001001001001;
				18'b010010000100100111: oled_data = 16'b1101010001010001;
				18'b010010000110100111: oled_data = 16'b1110110011110011;
				18'b010010001000100111: oled_data = 16'b1100001100001101;
				18'b010010001010100111: oled_data = 16'b1011001000101001;
				18'b010010001100100111: oled_data = 16'b1011001000101001;
				18'b010010001110100111: oled_data = 16'b1011001001001001;
				18'b010010010000100111: oled_data = 16'b1011001001101010;
				18'b010010010010100111: oled_data = 16'b1011001000101001;
				18'b010010010100100111: oled_data = 16'b1011101111110000;
				18'b010010010110100111: oled_data = 16'b1100011100011100;
				18'b010010011000100111: oled_data = 16'b1011110111010111;
				18'b010010011010100111: oled_data = 16'b1011001001001001;
				18'b010010011100100111: oled_data = 16'b1011001000101001;
				18'b010010011110100111: oled_data = 16'b1011001001001001;
				18'b010010100000100111: oled_data = 16'b1011001000101000;
				18'b010010100010100111: oled_data = 16'b1010101000001000;
				18'b010010100100100111: oled_data = 16'b1010000111101000;
				18'b010010100110100111: oled_data = 16'b1010101000001000;
				18'b010000011000101000: oled_data = 16'b0011000110100101;
				18'b010000011010101000: oled_data = 16'b0100101000100110;
				18'b010000011100101000: oled_data = 16'b0101101011001001;
				18'b010000011110101000: oled_data = 16'b0110101101001100;
				18'b010000100000101000: oled_data = 16'b1000101111110000;
				18'b010000100010101000: oled_data = 16'b1010101110010000;
				18'b010000100100101000: oled_data = 16'b1011001101010000;
				18'b010000100110101000: oled_data = 16'b1011001101110001;
				18'b010000101000101000: oled_data = 16'b1101110010110110;
				18'b010000101010101000: oled_data = 16'b1101110011010110;
				18'b010000101100101000: oled_data = 16'b1101110011010101;
				18'b010000101110101000: oled_data = 16'b1110011010011001;
				18'b010000110000101000: oled_data = 16'b1110011100011011;
				18'b010000110010101000: oled_data = 16'b1110011010111010;
				18'b010000110100101000: oled_data = 16'b1101010100010101;
				18'b010000110110101000: oled_data = 16'b1110010011010110;
				18'b010000111000101000: oled_data = 16'b1101110011010101;
				18'b010000111010101000: oled_data = 16'b1101110011010110;
				18'b010000111100101000: oled_data = 16'b1101110011010101;
				18'b010000111110101000: oled_data = 16'b1101110011010101;
				18'b010001000000101000: oled_data = 16'b1101110011010101;
				18'b010001000010101000: oled_data = 16'b1101110011010101;
				18'b010001000100101000: oled_data = 16'b1101110010110101;
				18'b010001000110101000: oled_data = 16'b1101010101010110;
				18'b010001001000101000: oled_data = 16'b1110111100011011;
				18'b010001001010101000: oled_data = 16'b1110111100011011;
				18'b010001001100101000: oled_data = 16'b1110111100011011;
				18'b010001001110101000: oled_data = 16'b1110111100011011;
				18'b010001010000101000: oled_data = 16'b1110011100011011;
				18'b010001010010101000: oled_data = 16'b1111011100111100;
				18'b010001010100101000: oled_data = 16'b1010110011110011;
				18'b010001010110101000: oled_data = 16'b0011100101000101;
				18'b010001011000101000: oled_data = 16'b0011100110000110;
				18'b010001011010101000: oled_data = 16'b1011010100110100;
				18'b010001011100101000: oled_data = 16'b1111011100111100;
				18'b010001011110101000: oled_data = 16'b1110111100011011;
				18'b010001100000101000: oled_data = 16'b1110111100011010;
				18'b010001100010101000: oled_data = 16'b1110111100011010;
				18'b010001100100101000: oled_data = 16'b1110111100011010;
				18'b010001100110101000: oled_data = 16'b1110111100011010;
				18'b010001101000101000: oled_data = 16'b1110111100011010;
				18'b010001101010101000: oled_data = 16'b1110111100011010;
				18'b010001101100101000: oled_data = 16'b1110111100011010;
				18'b010001101110101000: oled_data = 16'b1110111100011011;
				18'b010001110000101000: oled_data = 16'b1101111010111001;
				18'b010001110010101000: oled_data = 16'b1110011011111010;
				18'b010001110100101000: oled_data = 16'b1110111100011011;
				18'b010001110110101000: oled_data = 16'b1110011011011001;
				18'b010001111000101000: oled_data = 16'b1101010110110110;
				18'b010001111010101000: oled_data = 16'b1101010101010101;
				18'b010001111100101000: oled_data = 16'b1101110100010100;
				18'b010001111110101000: oled_data = 16'b1100101111001111;
				18'b010010000000101000: oled_data = 16'b1010101000001000;
				18'b010010000010101000: oled_data = 16'b1011101011101100;
				18'b010010000100101000: oled_data = 16'b1110110011110100;
				18'b010010000110101000: oled_data = 16'b1100101101101110;
				18'b010010001000101000: oled_data = 16'b1011001000101001;
				18'b010010001010101000: oled_data = 16'b1011001001001001;
				18'b010010001100101000: oled_data = 16'b1011001001001001;
				18'b010010001110101000: oled_data = 16'b1011001001001001;
				18'b010010010000101000: oled_data = 16'b1011001001001001;
				18'b010010010010101000: oled_data = 16'b1011001001001001;
				18'b010010010100101000: oled_data = 16'b1100010110110110;
				18'b010010010110101000: oled_data = 16'b1011111100011100;
				18'b010010011000101000: oled_data = 16'b1011111011111011;
				18'b010010011010101000: oled_data = 16'b1011001101101110;
				18'b010010011100101000: oled_data = 16'b1010101000001000;
				18'b010010011110101000: oled_data = 16'b1010101000001000;
				18'b010010100000101000: oled_data = 16'b1010001000001000;
				18'b010010100010101000: oled_data = 16'b1010001000001000;
				18'b010010100100101000: oled_data = 16'b1010101000001000;
				18'b010010100110101000: oled_data = 16'b1010101000001000;
				18'b010000011000101001: oled_data = 16'b0111001110001010;
				18'b010000011010101001: oled_data = 16'b0111101110101010;
				18'b010000011100101001: oled_data = 16'b0111101111101011;
				18'b010000011110101001: oled_data = 16'b0110101101001100;
				18'b010000100000101001: oled_data = 16'b0110101011001100;
				18'b010000100010101001: oled_data = 16'b1011001110010001;
				18'b010000100100101001: oled_data = 16'b1010101100110000;
				18'b010000100110101001: oled_data = 16'b1100110000110011;
				18'b010000101000101001: oled_data = 16'b1110010011010110;
				18'b010000101010101001: oled_data = 16'b1101110011010110;
				18'b010000101100101001: oled_data = 16'b1101110011010101;
				18'b010000101110101001: oled_data = 16'b1110011001111001;
				18'b010000110000101001: oled_data = 16'b1110111100011011;
				18'b010000110010101001: oled_data = 16'b1110011011011010;
				18'b010000110100101001: oled_data = 16'b1101010100010101;
				18'b010000110110101001: oled_data = 16'b1110010011010110;
				18'b010000111000101001: oled_data = 16'b1101110011010110;
				18'b010000111010101001: oled_data = 16'b1110010011010110;
				18'b010000111100101001: oled_data = 16'b1101110011010101;
				18'b010000111110101001: oled_data = 16'b1101110011010101;
				18'b010001000000101001: oled_data = 16'b1101110011010101;
				18'b010001000010101001: oled_data = 16'b1101110011010101;
				18'b010001000100101001: oled_data = 16'b1101110010110101;
				18'b010001000110101001: oled_data = 16'b1101010100110110;
				18'b010001001000101001: oled_data = 16'b1110011011111010;
				18'b010001001010101001: oled_data = 16'b1110111100011010;
				18'b010001001100101001: oled_data = 16'b1110111100011010;
				18'b010001001110101001: oled_data = 16'b1110111100011010;
				18'b010001010000101001: oled_data = 16'b1111011101011011;
				18'b010001010010101001: oled_data = 16'b1011010101010100;
				18'b010001010100101001: oled_data = 16'b0011100110000101;
				18'b010001010110101001: oled_data = 16'b0011100110000110;
				18'b010001011000101001: oled_data = 16'b1010110100110100;
				18'b010001011010101001: oled_data = 16'b1110111100111100;
				18'b010001011100101001: oled_data = 16'b1110111011111011;
				18'b010001011110101001: oled_data = 16'b1110111100011011;
				18'b010001100000101001: oled_data = 16'b1110111100011010;
				18'b010001100010101001: oled_data = 16'b1110111100011010;
				18'b010001100100101001: oled_data = 16'b1110011100011010;
				18'b010001100110101001: oled_data = 16'b1110111100011010;
				18'b010001101000101001: oled_data = 16'b1110111100011010;
				18'b010001101010101001: oled_data = 16'b1110111100011010;
				18'b010001101100101001: oled_data = 16'b1110111100011010;
				18'b010001101110101001: oled_data = 16'b1101111010111001;
				18'b010001110000101001: oled_data = 16'b1110011011011010;
				18'b010001110010101001: oled_data = 16'b1110111100111011;
				18'b010001110100101001: oled_data = 16'b1110011011011010;
				18'b010001110110101001: oled_data = 16'b1100010101010100;
				18'b010001111000101001: oled_data = 16'b1101010111110110;
				18'b010001111010101001: oled_data = 16'b1110011010011001;
				18'b010001111100101001: oled_data = 16'b1101110100010100;
				18'b010001111110101001: oled_data = 16'b1100101110001110;
				18'b010010000000101001: oled_data = 16'b1011001000001000;
				18'b010010000010101001: oled_data = 16'b1100101110101110;
				18'b010010000100101001: oled_data = 16'b1110010011010010;
				18'b010010000110101001: oled_data = 16'b1011101010001010;
				18'b010010001000101001: oled_data = 16'b1011001001001001;
				18'b010010001010101001: oled_data = 16'b1011001001001001;
				18'b010010001100101001: oled_data = 16'b1011001001001001;
				18'b010010001110101001: oled_data = 16'b1011001001001001;
				18'b010010010000101001: oled_data = 16'b1011001000101001;
				18'b010010010010101001: oled_data = 16'b1011001101101110;
				18'b010010010100101001: oled_data = 16'b1100011011011011;
				18'b010010010110101001: oled_data = 16'b1011111011111011;
				18'b010010011000101001: oled_data = 16'b1011111100011100;
				18'b010010011010101001: oled_data = 16'b1011110101010101;
				18'b010010011100101001: oled_data = 16'b1010101000101001;
				18'b010010011110101001: oled_data = 16'b1011001000101000;
				18'b010010100000101001: oled_data = 16'b1011001000101000;
				18'b010010100010101001: oled_data = 16'b1010101000101000;
				18'b010010100100101001: oled_data = 16'b1010101000001000;
				18'b010010100110101001: oled_data = 16'b1010101000001000;
				18'b010000011000101010: oled_data = 16'b0111101110101011;
				18'b010000011010101010: oled_data = 16'b0101101011001000;
				18'b010000011100101010: oled_data = 16'b0111001101101010;
				18'b010000011110101010: oled_data = 16'b0111001100101100;
				18'b010000100000101010: oled_data = 16'b1010001110110000;
				18'b010000100010101010: oled_data = 16'b1011001110010001;
				18'b010000100100101010: oled_data = 16'b1100001111110010;
				18'b010000100110101010: oled_data = 16'b1101110011010101;
				18'b010000101000101010: oled_data = 16'b1101110011010110;
				18'b010000101010101010: oled_data = 16'b1101110011010101;
				18'b010000101100101010: oled_data = 16'b1101110010110101;
				18'b010000101110101010: oled_data = 16'b1101010110110111;
				18'b010000110000101010: oled_data = 16'b1110111100011011;
				18'b010000110010101010: oled_data = 16'b1110011011011010;
				18'b010000110100101010: oled_data = 16'b1101010100010101;
				18'b010000110110101010: oled_data = 16'b1110010011010110;
				18'b010000111000101010: oled_data = 16'b1110010011010110;
				18'b010000111010101010: oled_data = 16'b1101110011010110;
				18'b010000111100101010: oled_data = 16'b1101110011010101;
				18'b010000111110101010: oled_data = 16'b1101110011010101;
				18'b010001000000101010: oled_data = 16'b1101110011010101;
				18'b010001000010101010: oled_data = 16'b1101110011010101;
				18'b010001000100101010: oled_data = 16'b1101110011010101;
				18'b010001000110101010: oled_data = 16'b1101010101010110;
				18'b010001001000101010: oled_data = 16'b1110011011111010;
				18'b010001001010101010: oled_data = 16'b1110111100011011;
				18'b010001001100101010: oled_data = 16'b1110111100011011;
				18'b010001001110101010: oled_data = 16'b1111011100111100;
				18'b010001010000101010: oled_data = 16'b1011010100110100;
				18'b010001010010101010: oled_data = 16'b0011100110000110;
				18'b010001010100101010: oled_data = 16'b0100000111000111;
				18'b010001010110101010: oled_data = 16'b1011010101110101;
				18'b010001011000101010: oled_data = 16'b1110111100111100;
				18'b010001011010101010: oled_data = 16'b1110111100011010;
				18'b010001011100101010: oled_data = 16'b1110111100011010;
				18'b010001011110101010: oled_data = 16'b1110111100011010;
				18'b010001100000101010: oled_data = 16'b1110111100011010;
				18'b010001100010101010: oled_data = 16'b1110111100011010;
				18'b010001100100101010: oled_data = 16'b1110111100011010;
				18'b010001100110101010: oled_data = 16'b1110111100011010;
				18'b010001101000101010: oled_data = 16'b1110111100011010;
				18'b010001101010101010: oled_data = 16'b1110111100011010;
				18'b010001101100101010: oled_data = 16'b1110111100011010;
				18'b010001101110101010: oled_data = 16'b1110011011111010;
				18'b010001110000101010: oled_data = 16'b1110111100111011;
				18'b010001110010101010: oled_data = 16'b1110011010111001;
				18'b010001110100101010: oled_data = 16'b1100110101010101;
				18'b010001110110101010: oled_data = 16'b1101010111110111;
				18'b010001111000101010: oled_data = 16'b1110011011111010;
				18'b010001111010101010: oled_data = 16'b1110011010111010;
				18'b010001111100101010: oled_data = 16'b1101010100010100;
				18'b010001111110101010: oled_data = 16'b1100001101001101;
				18'b010010000000101010: oled_data = 16'b1010101000101000;
				18'b010010000010101010: oled_data = 16'b1101010000110000;
				18'b010010000100101010: oled_data = 16'b1101110000010000;
				18'b010010000110101010: oled_data = 16'b1011001001001001;
				18'b010010001000101010: oled_data = 16'b1011101001001001;
				18'b010010001010101010: oled_data = 16'b1011001001001001;
				18'b010010001100101010: oled_data = 16'b1011001001001001;
				18'b010010001110101010: oled_data = 16'b1011001001001001;
				18'b010010010000101010: oled_data = 16'b1011001000101001;
				18'b010010010010101010: oled_data = 16'b1011110101110110;
				18'b010010010100101010: oled_data = 16'b1011111100011100;
				18'b010010010110101010: oled_data = 16'b1011111011111011;
				18'b010010011000101010: oled_data = 16'b1011111011111100;
				18'b010010011010101010: oled_data = 16'b1100011010111011;
				18'b010010011100101010: oled_data = 16'b1011001100001100;
				18'b010010011110101010: oled_data = 16'b1010101000101000;
				18'b010010100000101010: oled_data = 16'b1011001000101001;
				18'b010010100010101010: oled_data = 16'b1010101000101000;
				18'b010010100100101010: oled_data = 16'b1010101000001000;
				18'b010010100110101010: oled_data = 16'b1010101000001000;
				18'b010000011000101011: oled_data = 16'b0111101110101011;
				18'b010000011010101011: oled_data = 16'b0111001110001011;
				18'b010000011100101011: oled_data = 16'b1000010000001101;
				18'b010000011110101011: oled_data = 16'b1001110000010000;
				18'b010000100000101011: oled_data = 16'b1101110010110101;
				18'b010000100010101011: oled_data = 16'b1100110001010100;
				18'b010000100100101011: oled_data = 16'b1101110011010110;
				18'b010000100110101011: oled_data = 16'b1101110011010101;
				18'b010000101000101011: oled_data = 16'b1101110011010101;
				18'b010000101010101011: oled_data = 16'b1101110011010101;
				18'b010000101100101011: oled_data = 16'b1101110010110101;
				18'b010000101110101011: oled_data = 16'b1100010010010011;
				18'b010000110000101011: oled_data = 16'b1110111011111011;
				18'b010000110010101011: oled_data = 16'b1110011011011010;
				18'b010000110100101011: oled_data = 16'b1101010100010101;
				18'b010000110110101011: oled_data = 16'b1110010011010110;
				18'b010000111000101011: oled_data = 16'b1110010011010110;
				18'b010000111010101011: oled_data = 16'b1101110011010110;
				18'b010000111100101011: oled_data = 16'b1101110011010101;
				18'b010000111110101011: oled_data = 16'b1101110011010101;
				18'b010001000000101011: oled_data = 16'b1101110011010101;
				18'b010001000010101011: oled_data = 16'b1101110011010101;
				18'b010001000100101011: oled_data = 16'b1101110011010101;
				18'b010001000110101011: oled_data = 16'b1101010101010110;
				18'b010001001000101011: oled_data = 16'b1110011100011011;
				18'b010001001010101011: oled_data = 16'b1110111100011010;
				18'b010001001100101011: oled_data = 16'b1111011100111011;
				18'b010001001110101011: oled_data = 16'b1011110101110101;
				18'b010001010000101011: oled_data = 16'b0011100101000101;
				18'b010001010010101011: oled_data = 16'b0100101000001000;
				18'b010001010100101011: oled_data = 16'b1100010111010110;
				18'b010001010110101011: oled_data = 16'b1110111100111100;
				18'b010001011000101011: oled_data = 16'b1110111100011011;
				18'b010001011010101011: oled_data = 16'b1110111011111010;
				18'b010001011100101011: oled_data = 16'b1110111100011010;
				18'b010001011110101011: oled_data = 16'b1110111100011010;
				18'b010001100000101011: oled_data = 16'b1110111100011010;
				18'b010001100010101011: oled_data = 16'b1110111100011010;
				18'b010001100100101011: oled_data = 16'b1110111100011011;
				18'b010001100110101011: oled_data = 16'b1110111100011010;
				18'b010001101000101011: oled_data = 16'b1110111100011010;
				18'b010001101010101011: oled_data = 16'b1110111100011010;
				18'b010001101100101011: oled_data = 16'b1110111100011010;
				18'b010001101110101011: oled_data = 16'b1110111100011011;
				18'b010001110000101011: oled_data = 16'b1101111001011000;
				18'b010001110010101011: oled_data = 16'b1101010100110100;
				18'b010001110100101011: oled_data = 16'b1101110110010110;
				18'b010001110110101011: oled_data = 16'b1110011010111001;
				18'b010001111000101011: oled_data = 16'b1110111100011010;
				18'b010001111010101011: oled_data = 16'b1110011011011010;
				18'b010001111100101011: oled_data = 16'b1101110101010101;
				18'b010001111110101011: oled_data = 16'b1011101100001100;
				18'b010010000000101011: oled_data = 16'b1010101000101001;
				18'b010010000010101011: oled_data = 16'b1101110001110001;
				18'b010010000100101011: oled_data = 16'b1100101101101110;
				18'b010010000110101011: oled_data = 16'b1011001000101001;
				18'b010010001000101011: oled_data = 16'b1011101001001001;
				18'b010010001010101011: oled_data = 16'b1011001001001001;
				18'b010010001100101011: oled_data = 16'b1011001001001001;
				18'b010010001110101011: oled_data = 16'b1011001000101001;
				18'b010010010000101011: oled_data = 16'b1010101011001011;
				18'b010010010010101011: oled_data = 16'b1011111010111010;
				18'b010010010100101011: oled_data = 16'b1011111011111100;
				18'b010010010110101011: oled_data = 16'b1011111011111011;
				18'b010010011000101011: oled_data = 16'b1011111011111100;
				18'b010010011010101011: oled_data = 16'b1100011100111100;
				18'b010010011100101011: oled_data = 16'b1011110011010010;
				18'b010010011110101011: oled_data = 16'b1010101000001000;
				18'b010010100000101011: oled_data = 16'b1010101000101000;
				18'b010010100010101011: oled_data = 16'b1010101000001000;
				18'b010010100100101011: oled_data = 16'b1010101000001000;
				18'b010010100110101011: oled_data = 16'b1010101000001000;
				18'b010000011000101100: oled_data = 16'b1001010001001110;
				18'b010000011010101100: oled_data = 16'b1000010000101110;
				18'b010000011100101100: oled_data = 16'b1000001111101110;
				18'b010000011110101100: oled_data = 16'b1100010010010011;
				18'b010000100000101100: oled_data = 16'b1101010010010100;
				18'b010000100010101100: oled_data = 16'b1101110011010110;
				18'b010000100100101100: oled_data = 16'b1101110011010110;
				18'b010000100110101100: oled_data = 16'b1101110011010101;
				18'b010000101000101100: oled_data = 16'b1101110011010101;
				18'b010000101010101100: oled_data = 16'b1101110011010110;
				18'b010000101100101100: oled_data = 16'b1101010010010101;
				18'b010000101110101100: oled_data = 16'b1011001110010001;
				18'b010000110000101100: oled_data = 16'b1101010101010110;
				18'b010000110010101100: oled_data = 16'b1110111100011010;
				18'b010000110100101100: oled_data = 16'b1101010100010101;
				18'b010000110110101100: oled_data = 16'b1101110010110110;
				18'b010000111000101100: oled_data = 16'b1101110011010110;
				18'b010000111010101100: oled_data = 16'b1101110011010101;
				18'b010000111100101100: oled_data = 16'b1101110011010101;
				18'b010000111110101100: oled_data = 16'b1101110011010101;
				18'b010001000000101100: oled_data = 16'b1101110011010101;
				18'b010001000010101100: oled_data = 16'b1101110011010101;
				18'b010001000100101100: oled_data = 16'b1101110010110101;
				18'b010001000110101100: oled_data = 16'b1101010101010110;
				18'b010001001000101100: oled_data = 16'b1110011011111010;
				18'b010001001010101100: oled_data = 16'b1110111100011010;
				18'b010001001100101100: oled_data = 16'b1110011011011001;
				18'b010001001110101100: oled_data = 16'b0101001001001000;
				18'b010001010000101100: oled_data = 16'b0110001010101010;
				18'b010001010010101100: oled_data = 16'b1101011001111000;
				18'b010001010100101100: oled_data = 16'b1110111100111011;
				18'b010001010110101100: oled_data = 16'b1110111100011010;
				18'b010001011000101100: oled_data = 16'b1110111100011010;
				18'b010001011010101100: oled_data = 16'b1110111100011010;
				18'b010001011100101100: oled_data = 16'b1110111100011010;
				18'b010001011110101100: oled_data = 16'b1110111100011010;
				18'b010001100000101100: oled_data = 16'b1110111100011010;
				18'b010001100010101100: oled_data = 16'b1110111100011010;
				18'b010001100100101100: oled_data = 16'b1110111100011011;
				18'b010001100110101100: oled_data = 16'b1110011100011010;
				18'b010001101000101100: oled_data = 16'b1110011100011010;
				18'b010001101010101100: oled_data = 16'b1110111100111011;
				18'b010001101100101100: oled_data = 16'b1110011011011010;
				18'b010001101110101100: oled_data = 16'b1101010101110101;
				18'b010001110000101100: oled_data = 16'b1101010100110101;
				18'b010001110010101100: oled_data = 16'b1101110101010101;
				18'b010001110100101100: oled_data = 16'b1101111000111000;
				18'b010001110110101100: oled_data = 16'b1110111100011010;
				18'b010001111000101100: oled_data = 16'b1110011100011010;
				18'b010001111010101100: oled_data = 16'b1110011100011010;
				18'b010001111100101100: oled_data = 16'b1101110101110101;
				18'b010001111110101100: oled_data = 16'b1011101011101100;
				18'b010010000000101100: oled_data = 16'b1011001001001001;
				18'b010010000010101100: oled_data = 16'b1101110010010010;
				18'b010010000100101100: oled_data = 16'b1100001011101100;
				18'b010010000110101100: oled_data = 16'b1011001000101001;
				18'b010010001000101100: oled_data = 16'b1011001001001001;
				18'b010010001010101100: oled_data = 16'b1011001001001001;
				18'b010010001100101100: oled_data = 16'b1011001001001001;
				18'b010010001110101100: oled_data = 16'b1011001000101001;
				18'b010010010000101100: oled_data = 16'b1011110000110001;
				18'b010010010010101100: oled_data = 16'b1100011100011100;
				18'b010010010100101100: oled_data = 16'b1011111011111011;
				18'b010010010110101100: oled_data = 16'b1011111011111011;
				18'b010010011000101100: oled_data = 16'b1011111011111100;
				18'b010010011010101100: oled_data = 16'b1100111100111101;
				18'b010010011100101100: oled_data = 16'b1011111000111000;
				18'b010010011110101100: oled_data = 16'b1010101010001010;
				18'b010010100000101100: oled_data = 16'b1010101000101000;
				18'b010010100010101100: oled_data = 16'b1010101000001000;
				18'b010010100100101100: oled_data = 16'b1010101000001000;
				18'b010010100110101100: oled_data = 16'b1010101000001000;
				18'b010000011000101101: oled_data = 16'b0110101100001010;
				18'b010000011010101101: oled_data = 16'b0100001001000111;
				18'b010000011100101101: oled_data = 16'b1000001101001110;
				18'b010000011110101101: oled_data = 16'b1101010011010101;
				18'b010000100000101101: oled_data = 16'b1101110010110101;
				18'b010000100010101101: oled_data = 16'b1101110011010101;
				18'b010000100100101101: oled_data = 16'b1101110011010110;
				18'b010000100110101101: oled_data = 16'b1101110011010101;
				18'b010000101000101101: oled_data = 16'b1101110011010101;
				18'b010000101010101101: oled_data = 16'b1101110011010110;
				18'b010000101100101101: oled_data = 16'b1101010001010100;
				18'b010000101110101101: oled_data = 16'b1011001101010000;
				18'b010000110000101101: oled_data = 16'b1011001110110001;
				18'b010000110010101101: oled_data = 16'b1101010111010111;
				18'b010000110100101101: oled_data = 16'b1101010011010101;
				18'b010000110110101101: oled_data = 16'b1101110010110110;
				18'b010000111000101101: oled_data = 16'b1101110011010101;
				18'b010000111010101101: oled_data = 16'b1101110011010101;
				18'b010000111100101101: oled_data = 16'b1101110011010101;
				18'b010000111110101101: oled_data = 16'b1101110011010101;
				18'b010001000000101101: oled_data = 16'b1101110011010101;
				18'b010001000010101101: oled_data = 16'b1101110011010101;
				18'b010001000100101101: oled_data = 16'b1101110010110101;
				18'b010001000110101101: oled_data = 16'b1101010101010110;
				18'b010001001000101101: oled_data = 16'b1110011011111010;
				18'b010001001010101101: oled_data = 16'b1110111100111011;
				18'b010001001100101101: oled_data = 16'b1011110110010100;
				18'b010001001110101101: oled_data = 16'b1000001110101101;
				18'b010001010000101101: oled_data = 16'b1110011011011010;
				18'b010001010010101101: oled_data = 16'b1110111100111011;
				18'b010001010100101101: oled_data = 16'b1110111100011010;
				18'b010001010110101101: oled_data = 16'b1110111100011010;
				18'b010001011000101101: oled_data = 16'b1110111100011010;
				18'b010001011010101101: oled_data = 16'b1110111100011010;
				18'b010001011100101101: oled_data = 16'b1110111100011010;
				18'b010001011110101101: oled_data = 16'b1110111100011010;
				18'b010001100000101101: oled_data = 16'b1110111100011010;
				18'b010001100010101101: oled_data = 16'b1110111100011010;
				18'b010001100100101101: oled_data = 16'b1110111100011010;
				18'b010001100110101101: oled_data = 16'b1110111100011010;
				18'b010001101000101101: oled_data = 16'b1110111100011010;
				18'b010001101010101101: oled_data = 16'b1101111000010111;
				18'b010001101100101101: oled_data = 16'b1011110001010001;
				18'b010001101110101101: oled_data = 16'b1100110010110011;
				18'b010001110000101101: oled_data = 16'b1110010101010101;
				18'b010001110010101101: oled_data = 16'b1101110100110101;
				18'b010001110100101101: oled_data = 16'b1110011001111000;
				18'b010001110110101101: oled_data = 16'b1110111100011010;
				18'b010001111000101101: oled_data = 16'b1110011100011010;
				18'b010001111010101101: oled_data = 16'b1110111100011011;
				18'b010001111100101101: oled_data = 16'b1101010110110110;
				18'b010001111110101101: oled_data = 16'b1011101011001100;
				18'b010010000000101101: oled_data = 16'b1011101001001010;
				18'b010010000010101101: oled_data = 16'b1101110001110001;
				18'b010010000100101101: oled_data = 16'b1011101010101011;
				18'b010010000110101101: oled_data = 16'b1011001001001001;
				18'b010010001000101101: oled_data = 16'b1011001001001001;
				18'b010010001010101101: oled_data = 16'b1011001001001001;
				18'b010010001100101101: oled_data = 16'b1011001001001001;
				18'b010010001110101101: oled_data = 16'b1011001001001001;
				18'b010010010000101101: oled_data = 16'b1100010110010111;
				18'b010010010010101101: oled_data = 16'b1011111100011100;
				18'b010010010100101101: oled_data = 16'b1011111011111011;
				18'b010010010110101101: oled_data = 16'b1011111011111011;
				18'b010010011000101101: oled_data = 16'b1011111011111100;
				18'b010010011010101101: oled_data = 16'b1100111100011101;
				18'b010010011100101101: oled_data = 16'b1011111011111011;
				18'b010010011110101101: oled_data = 16'b1010101101101101;
				18'b010010100000101101: oled_data = 16'b1010101000001000;
				18'b010010100010101101: oled_data = 16'b1010101000001000;
				18'b010010100100101101: oled_data = 16'b1010101000001000;
				18'b010010100110101101: oled_data = 16'b1010101000001000;
				18'b010000011000101110: oled_data = 16'b0100000111100111;
				18'b010000011010101110: oled_data = 16'b0110101010101011;
				18'b010000011100101110: oled_data = 16'b1100110001110100;
				18'b010000011110101110: oled_data = 16'b1101110010010101;
				18'b010000100000101110: oled_data = 16'b1101110010110101;
				18'b010000100010101110: oled_data = 16'b1101110010110101;
				18'b010000100100101110: oled_data = 16'b1101110010110101;
				18'b010000100110101110: oled_data = 16'b1101110010110101;
				18'b010000101000101110: oled_data = 16'b1101110010110101;
				18'b010000101010101110: oled_data = 16'b1101110011010101;
				18'b010000101100101110: oled_data = 16'b1100001111110010;
				18'b010000101110101110: oled_data = 16'b1011001101010000;
				18'b010000110000101110: oled_data = 16'b1011001101010000;
				18'b010000110010101110: oled_data = 16'b1010101101110000;
				18'b010000110100101110: oled_data = 16'b1100110001110100;
				18'b010000110110101110: oled_data = 16'b1101110011010101;
				18'b010000111000101110: oled_data = 16'b1101110010110101;
				18'b010000111010101110: oled_data = 16'b1101110010110110;
				18'b010000111100101110: oled_data = 16'b1101110011010101;
				18'b010000111110101110: oled_data = 16'b1101110011010101;
				18'b010001000000101110: oled_data = 16'b1101110010110101;
				18'b010001000010101110: oled_data = 16'b1101110010110101;
				18'b010001000100101110: oled_data = 16'b1101110010110101;
				18'b010001000110101110: oled_data = 16'b1101110101010110;
				18'b010001001000101110: oled_data = 16'b1110011100011010;
				18'b010001001010101110: oled_data = 16'b1110011100011010;
				18'b010001001100101110: oled_data = 16'b1110011011011001;
				18'b010001001110101110: oled_data = 16'b1110011100011010;
				18'b010001010000101110: oled_data = 16'b1110111100011011;
				18'b010001010010101110: oled_data = 16'b1110111100011010;
				18'b010001010100101110: oled_data = 16'b1110111100011010;
				18'b010001010110101110: oled_data = 16'b1110011100011010;
				18'b010001011000101110: oled_data = 16'b1110011100011011;
				18'b010001011010101110: oled_data = 16'b1110011100011010;
				18'b010001011100101110: oled_data = 16'b1110011100011010;
				18'b010001011110101110: oled_data = 16'b1110111100011010;
				18'b010001100000101110: oled_data = 16'b1110111100011010;
				18'b010001100010101110: oled_data = 16'b1110111100011010;
				18'b010001100100101110: oled_data = 16'b1110111100011010;
				18'b010001100110101110: oled_data = 16'b1101111000110111;
				18'b010001101000101110: oled_data = 16'b1100010011010011;
				18'b010001101010101110: oled_data = 16'b1011001110001111;
				18'b010001101100101110: oled_data = 16'b1100001111110001;
				18'b010001101110101110: oled_data = 16'b1101110100010101;
				18'b010001110000101110: oled_data = 16'b1101110101010101;
				18'b010001110010101110: oled_data = 16'b1101110101010101;
				18'b010001110100101110: oled_data = 16'b1110011010011001;
				18'b010001110110101110: oled_data = 16'b1110111100011010;
				18'b010001111000101110: oled_data = 16'b1110011100011010;
				18'b010001111010101110: oled_data = 16'b1110111100011010;
				18'b010001111100101110: oled_data = 16'b1101111000110111;
				18'b010001111110101110: oled_data = 16'b1011001011001011;
				18'b010010000000101110: oled_data = 16'b1011001001101010;
				18'b010010000010101110: oled_data = 16'b1101010000110000;
				18'b010010000100101110: oled_data = 16'b1011101001101010;
				18'b010010000110101110: oled_data = 16'b1011001001001001;
				18'b010010001000101110: oled_data = 16'b1011001001001001;
				18'b010010001010101110: oled_data = 16'b1011001001001001;
				18'b010010001100101110: oled_data = 16'b1011001000101001;
				18'b010010001110101110: oled_data = 16'b1011001010001010;
				18'b010010010000101110: oled_data = 16'b1100011001011001;
				18'b010010010010101110: oled_data = 16'b1011111011111100;
				18'b010010010100101110: oled_data = 16'b1011111011011011;
				18'b010010010110101110: oled_data = 16'b1011111011011011;
				18'b010010011000101110: oled_data = 16'b1011111011011011;
				18'b010010011010101110: oled_data = 16'b1100111100011100;
				18'b010010011100101110: oled_data = 16'b1011111100011100;
				18'b010010011110101110: oled_data = 16'b1011010010010010;
				18'b010010100000101110: oled_data = 16'b1010100111101000;
				18'b010010100010101110: oled_data = 16'b1010101000001000;
				18'b010010100100101110: oled_data = 16'b1010101000001000;
				18'b010010100110101110: oled_data = 16'b1010101000001000;
				18'b010000011000101111: oled_data = 16'b0110001001101001;
				18'b010000011010101111: oled_data = 16'b1011110000010010;
				18'b010000011100101111: oled_data = 16'b1101010010010101;
				18'b010000011110101111: oled_data = 16'b1101110010110101;
				18'b010000100000101111: oled_data = 16'b1101110010110101;
				18'b010000100010101111: oled_data = 16'b1101110010110101;
				18'b010000100100101111: oled_data = 16'b1101110010010101;
				18'b010000100110101111: oled_data = 16'b1101110010010101;
				18'b010000101000101111: oled_data = 16'b1101110010110101;
				18'b010000101010101111: oled_data = 16'b1101110010110101;
				18'b010000101100101111: oled_data = 16'b1011101110110001;
				18'b010000101110101111: oled_data = 16'b1011001101010000;
				18'b010000110000101111: oled_data = 16'b1011001101110000;
				18'b010000110010101111: oled_data = 16'b1011001101010000;
				18'b010000110100101111: oled_data = 16'b1101010001010100;
				18'b010000110110101111: oled_data = 16'b1101110010110101;
				18'b010000111000101111: oled_data = 16'b1101110010110101;
				18'b010000111010101111: oled_data = 16'b1101110010110101;
				18'b010000111100101111: oled_data = 16'b1101110010110101;
				18'b010000111110101111: oled_data = 16'b1101110010110101;
				18'b010001000000101111: oled_data = 16'b1101110010110101;
				18'b010001000010101111: oled_data = 16'b1101110010110101;
				18'b010001000100101111: oled_data = 16'b1101110010010101;
				18'b010001000110101111: oled_data = 16'b1101110110010111;
				18'b010001001000101111: oled_data = 16'b1110011011111010;
				18'b010001001010101111: oled_data = 16'b1110011011111010;
				18'b010001001100101111: oled_data = 16'b1110011011111010;
				18'b010001001110101111: oled_data = 16'b1110111100011010;
				18'b010001010000101111: oled_data = 16'b1110011100011010;
				18'b010001010010101111: oled_data = 16'b1110011011111010;
				18'b010001010100101111: oled_data = 16'b1110011011111010;
				18'b010001010110101111: oled_data = 16'b1110011011111010;
				18'b010001011000101111: oled_data = 16'b1110011011111010;
				18'b010001011010101111: oled_data = 16'b1110011100011010;
				18'b010001011100101111: oled_data = 16'b1110111100011010;
				18'b010001011110101111: oled_data = 16'b1110111100011010;
				18'b010001100000101111: oled_data = 16'b1110011010111001;
				18'b010001100010101111: oled_data = 16'b1101010111010110;
				18'b010001100100101111: oled_data = 16'b1011110010110010;
				18'b010001100110101111: oled_data = 16'b1011001110101111;
				18'b010001101000101111: oled_data = 16'b1011101110001111;
				18'b010001101010101111: oled_data = 16'b1011001110101111;
				18'b010001101100101111: oled_data = 16'b1101010011010100;
				18'b010001101110101111: oled_data = 16'b1110010100110101;
				18'b010001110000101111: oled_data = 16'b1101110100110101;
				18'b010001110010101111: oled_data = 16'b1101010101110110;
				18'b010001110100101111: oled_data = 16'b1110011011011010;
				18'b010001110110101111: oled_data = 16'b1110111100011010;
				18'b010001111000101111: oled_data = 16'b1110011011111010;
				18'b010001111010101111: oled_data = 16'b1110011100011010;
				18'b010001111100101111: oled_data = 16'b1110011011111001;
				18'b010001111110101111: oled_data = 16'b1010101100101100;
				18'b010010000000101111: oled_data = 16'b1011001001101010;
				18'b010010000010101111: oled_data = 16'b1100101111101111;
				18'b010010000100101111: oled_data = 16'b1011001001001001;
				18'b010010000110101111: oled_data = 16'b1011001001001001;
				18'b010010001000101111: oled_data = 16'b1011001001101001;
				18'b010010001010101111: oled_data = 16'b1011001001001001;
				18'b010010001100101111: oled_data = 16'b1011001000101000;
				18'b010010001110101111: oled_data = 16'b1011101011101100;
				18'b010010010000101111: oled_data = 16'b1100011010111011;
				18'b010010010010101111: oled_data = 16'b1011111011011100;
				18'b010010010100101111: oled_data = 16'b1011111011011011;
				18'b010010010110101111: oled_data = 16'b1011111011011011;
				18'b010010011000101111: oled_data = 16'b1011111011011100;
				18'b010010011010101111: oled_data = 16'b1100011011111100;
				18'b010010011100101111: oled_data = 16'b1011111100011100;
				18'b010010011110101111: oled_data = 16'b1011110100010100;
				18'b010010100000101111: oled_data = 16'b1010100111101000;
				18'b010010100010101111: oled_data = 16'b1010100111101000;
				18'b010010100100101111: oled_data = 16'b1010101000001000;
				18'b010010100110101111: oled_data = 16'b1010100111101000;
				18'b010000011000110000: oled_data = 16'b1010101111010001;
				18'b010000011010110000: oled_data = 16'b1100110001010100;
				18'b010000011100110000: oled_data = 16'b1101110010110101;
				18'b010000011110110000: oled_data = 16'b1101110010010101;
				18'b010000100000110000: oled_data = 16'b1101110010010101;
				18'b010000100010110000: oled_data = 16'b1101010010010101;
				18'b010000100100110000: oled_data = 16'b1101010010010101;
				18'b010000100110110000: oled_data = 16'b1101010010010101;
				18'b010000101000110000: oled_data = 16'b1101110010010101;
				18'b010000101010110000: oled_data = 16'b1100110000110011;
				18'b010000101100110000: oled_data = 16'b1010101100101111;
				18'b010000101110110000: oled_data = 16'b1011001101010000;
				18'b010000110000110000: oled_data = 16'b1011001101010000;
				18'b010000110010110000: oled_data = 16'b1010101100110000;
				18'b010000110100110000: oled_data = 16'b1101010001010100;
				18'b010000110110110000: oled_data = 16'b1101110010010101;
				18'b010000111000110000: oled_data = 16'b1101010010010101;
				18'b010000111010110000: oled_data = 16'b1101110010010101;
				18'b010000111100110000: oled_data = 16'b1101110010110101;
				18'b010000111110110000: oled_data = 16'b1101110010110101;
				18'b010001000000110000: oled_data = 16'b1101110010110101;
				18'b010001000010110000: oled_data = 16'b1101110010110101;
				18'b010001000100110000: oled_data = 16'b1101010010010101;
				18'b010001000110110000: oled_data = 16'b1101110111011000;
				18'b010001001000110000: oled_data = 16'b1110011100011010;
				18'b010001001010110000: oled_data = 16'b1110011100011010;
				18'b010001001100110000: oled_data = 16'b1110011011111010;
				18'b010001001110110000: oled_data = 16'b1110011011011010;
				18'b010001010000110000: oled_data = 16'b1110011011011010;
				18'b010001010010110000: oled_data = 16'b1110011011011010;
				18'b010001010100110000: oled_data = 16'b1110011011111010;
				18'b010001010110110000: oled_data = 16'b1110011011111010;
				18'b010001011000110000: oled_data = 16'b1101111010111001;
				18'b010001011010110000: oled_data = 16'b1100110111110110;
				18'b010001011100110000: oled_data = 16'b1100110101110101;
				18'b010001011110110000: oled_data = 16'b1011110010110010;
				18'b010001100000110000: oled_data = 16'b1011001111110000;
				18'b010001100010110000: oled_data = 16'b1011001110001111;
				18'b010001100100110000: oled_data = 16'b1011001110001111;
				18'b010001100110110000: oled_data = 16'b1011101111010000;
				18'b010001101000110000: oled_data = 16'b1011001110001111;
				18'b010001101010110000: oled_data = 16'b1100110001010010;
				18'b010001101100110000: oled_data = 16'b1101110100110101;
				18'b010001101110110000: oled_data = 16'b1101110100110101;
				18'b010001110000110000: oled_data = 16'b1101110100010101;
				18'b010001110010110000: oled_data = 16'b1101010101110110;
				18'b010001110100110000: oled_data = 16'b1110011011011010;
				18'b010001110110110000: oled_data = 16'b1110111011111010;
				18'b010001111000110000: oled_data = 16'b1110011011111010;
				18'b010001111010110000: oled_data = 16'b1110011011111010;
				18'b010001111100110000: oled_data = 16'b1110011011111010;
				18'b010001111110110000: oled_data = 16'b1011001110101110;
				18'b010010000000110000: oled_data = 16'b1011001001101010;
				18'b010010000010110000: oled_data = 16'b1100101110001110;
				18'b010010000100110000: oled_data = 16'b1011001000101001;
				18'b010010000110110000: oled_data = 16'b1011001000101001;
				18'b010010001000110000: oled_data = 16'b1100101101101101;
				18'b010010001010110000: oled_data = 16'b1011101001101010;
				18'b010010001100110000: oled_data = 16'b1011001000101000;
				18'b010010001110110000: oled_data = 16'b1011101100001100;
				18'b010010010000110000: oled_data = 16'b1100011010111011;
				18'b010010010010110000: oled_data = 16'b1011111011011100;
				18'b010010010100110000: oled_data = 16'b1011111011011100;
				18'b010010010110110000: oled_data = 16'b1011011010111011;
				18'b010010011000110000: oled_data = 16'b1010111001111010;
				18'b010010011010110000: oled_data = 16'b1011011010111011;
				18'b010010011100110000: oled_data = 16'b1011111100011100;
				18'b010010011110110000: oled_data = 16'b1011110100110101;
				18'b010010100000110000: oled_data = 16'b1010100111001000;
				18'b010010100010110000: oled_data = 16'b1001100111000111;
				18'b010010100100110000: oled_data = 16'b1001100111000111;
				18'b010010100110110000: oled_data = 16'b1001100111000111;
				18'b010000011000110001: oled_data = 16'b1100110000110011;
				18'b010000011010110001: oled_data = 16'b1101010001110100;
				18'b010000011100110001: oled_data = 16'b1101010001110100;
				18'b010000011110110001: oled_data = 16'b1101010001110100;
				18'b010000100000110001: oled_data = 16'b1101010001110100;
				18'b010000100010110001: oled_data = 16'b1101010001110100;
				18'b010000100100110001: oled_data = 16'b1101010001110100;
				18'b010000100110110001: oled_data = 16'b1101010001110100;
				18'b010000101000110001: oled_data = 16'b1101010010010101;
				18'b010000101010110001: oled_data = 16'b1011101110010001;
				18'b010000101100110001: oled_data = 16'b1010101100101111;
				18'b010000101110110001: oled_data = 16'b1010101100010000;
				18'b010000110000110001: oled_data = 16'b1010101100001111;
				18'b010000110010110001: oled_data = 16'b1011001101110001;
				18'b010000110100110001: oled_data = 16'b1101010001110101;
				18'b010000110110110001: oled_data = 16'b1101010001110101;
				18'b010000111000110001: oled_data = 16'b1101010001110100;
				18'b010000111010110001: oled_data = 16'b1101010001110100;
				18'b010000111100110001: oled_data = 16'b1101010010010100;
				18'b010000111110110001: oled_data = 16'b1101010010010100;
				18'b010001000000110001: oled_data = 16'b1101010010010100;
				18'b010001000010110001: oled_data = 16'b1101010010010100;
				18'b010001000100110001: oled_data = 16'b1101010001110100;
				18'b010001000110110001: oled_data = 16'b1100110100110110;
				18'b010001001000110001: oled_data = 16'b1101010111110111;
				18'b010001001010110001: oled_data = 16'b1100110110110110;
				18'b010001001100110001: oled_data = 16'b1100110111110110;
				18'b010001001110110001: oled_data = 16'b1110011010111001;
				18'b010001010000110001: oled_data = 16'b1110011010111001;
				18'b010001010010110001: oled_data = 16'b1110011011011001;
				18'b010001010100110001: oled_data = 16'b1110011011111010;
				18'b010001010110110001: oled_data = 16'b1110011011111001;
				18'b010001011000110001: oled_data = 16'b1101111010111001;
				18'b010001011010110001: oled_data = 16'b1100110110110110;
				18'b010001011100110001: oled_data = 16'b1011010000010000;
				18'b010001011110110001: oled_data = 16'b1011001110001111;
				18'b010001100000110001: oled_data = 16'b1011101110110000;
				18'b010001100010110001: oled_data = 16'b1011001110001111;
				18'b010001100100110001: oled_data = 16'b1011001110010000;
				18'b010001100110110001: oled_data = 16'b1011101111010000;
				18'b010001101000110001: oled_data = 16'b1100010000010001;
				18'b010001101010110001: oled_data = 16'b1101110100010100;
				18'b010001101100110001: oled_data = 16'b1101110100010100;
				18'b010001101110110001: oled_data = 16'b1101110100010100;
				18'b010001110000110001: oled_data = 16'b1101110011110100;
				18'b010001110010110001: oled_data = 16'b1101010101110110;
				18'b010001110100110001: oled_data = 16'b1110011011011001;
				18'b010001110110110001: oled_data = 16'b1110011011011010;
				18'b010001111000110001: oled_data = 16'b1110011011111010;
				18'b010001111010110001: oled_data = 16'b1110011011011010;
				18'b010001111100110001: oled_data = 16'b1110011011011010;
				18'b010001111110110001: oled_data = 16'b1011001111001110;
				18'b010010000000110001: oled_data = 16'b1011001001101001;
				18'b010010000010110001: oled_data = 16'b1100001101001101;
				18'b010010000100110001: oled_data = 16'b1011001000101001;
				18'b010010000110110001: oled_data = 16'b1011001001001001;
				18'b010010001000110001: oled_data = 16'b1100101101101101;
				18'b010010001010110001: oled_data = 16'b1011001001001001;
				18'b010010001100110001: oled_data = 16'b1011001000001000;
				18'b010010001110110001: oled_data = 16'b1011101011101100;
				18'b010010010000110001: oled_data = 16'b1100011010111011;
				18'b010010010010110001: oled_data = 16'b1011111011111100;
				18'b010010010100110001: oled_data = 16'b1011011011011011;
				18'b010010010110110001: oled_data = 16'b1001110111111000;
				18'b010010011000110001: oled_data = 16'b1001010110111000;
				18'b010010011010110001: oled_data = 16'b1010111001111010;
				18'b010010011100110001: oled_data = 16'b1011111100011100;
				18'b010010011110110001: oled_data = 16'b1011010010010010;
				18'b010010100000110001: oled_data = 16'b1010000111000111;
				18'b010010100010110001: oled_data = 16'b1010000111101000;
				18'b010010100100110001: oled_data = 16'b1010000111100111;
				18'b010010100110110001: oled_data = 16'b1010000111000111;
				18'b010000011000110010: oled_data = 16'b1100110001010100;
				18'b010000011010110010: oled_data = 16'b1100110001010011;
				18'b010000011100110010: oled_data = 16'b1100110001010011;
				18'b010000011110110010: oled_data = 16'b1100110001010100;
				18'b010000100000110010: oled_data = 16'b1100110001010100;
				18'b010000100010110010: oled_data = 16'b1101010001010100;
				18'b010000100100110010: oled_data = 16'b1100110001010100;
				18'b010000100110110010: oled_data = 16'b1100110000110100;
				18'b010000101000110010: oled_data = 16'b1100110001010100;
				18'b010000101010110010: oled_data = 16'b1010101100001111;
				18'b010000101100110010: oled_data = 16'b1010101100001111;
				18'b010000101110110010: oled_data = 16'b1010101100001111;
				18'b010000110000110010: oled_data = 16'b1010001011101111;
				18'b010000110010110010: oled_data = 16'b1100001111110010;
				18'b010000110100110010: oled_data = 16'b1101010001110101;
				18'b010000110110110010: oled_data = 16'b1101010001110101;
				18'b010000111000110010: oled_data = 16'b1101010001110100;
				18'b010000111010110010: oled_data = 16'b1101010001110100;
				18'b010000111100110010: oled_data = 16'b1101010001110100;
				18'b010000111110110010: oled_data = 16'b1101010001110100;
				18'b010001000000110010: oled_data = 16'b1101010001110100;
				18'b010001000010110010: oled_data = 16'b1101010001110100;
				18'b010001000100110010: oled_data = 16'b1100110001010011;
				18'b010001000110110010: oled_data = 16'b1100010001010011;
				18'b010001001000110010: oled_data = 16'b1100010001010010;
				18'b010001001010110010: oled_data = 16'b1100010001110010;
				18'b010001001100110010: oled_data = 16'b1101011000010111;
				18'b010001001110110010: oled_data = 16'b1101111011011001;
				18'b010001010000110010: oled_data = 16'b1101111010111001;
				18'b010001010010110010: oled_data = 16'b1110011010111001;
				18'b010001010100110010: oled_data = 16'b1110011011011001;
				18'b010001010110110010: oled_data = 16'b1101111011011001;
				18'b010001011000110010: oled_data = 16'b1110011011011001;
				18'b010001011010110010: oled_data = 16'b1110011010111001;
				18'b010001011100110010: oled_data = 16'b1100110101010100;
				18'b010001011110110010: oled_data = 16'b1011001111110000;
				18'b010001100000110010: oled_data = 16'b1011101110110000;
				18'b010001100010110010: oled_data = 16'b1011001110001111;
				18'b010001100100110010: oled_data = 16'b1011101111110001;
				18'b010001100110110010: oled_data = 16'b1100010001010010;
				18'b010001101000110010: oled_data = 16'b1101010011110100;
				18'b010001101010110010: oled_data = 16'b1101110100010101;
				18'b010001101100110010: oled_data = 16'b1101010011110100;
				18'b010001101110110010: oled_data = 16'b1101010011110100;
				18'b010001110000110010: oled_data = 16'b1101010011010100;
				18'b010001110010110010: oled_data = 16'b1101110101110110;
				18'b010001110100110010: oled_data = 16'b1110011010111001;
				18'b010001110110110010: oled_data = 16'b1110011011011010;
				18'b010001111000110010: oled_data = 16'b1110011011011001;
				18'b010001111010110010: oled_data = 16'b1110011011011001;
				18'b010001111100110010: oled_data = 16'b1110011011011001;
				18'b010001111110110010: oled_data = 16'b1011001111001110;
				18'b010010000000110010: oled_data = 16'b1011001001001001;
				18'b010010000010110010: oled_data = 16'b1100001100101100;
				18'b010010000100110010: oled_data = 16'b1011001000101001;
				18'b010010000110110010: oled_data = 16'b1011001001001001;
				18'b010010001000110010: oled_data = 16'b1011101010101010;
				18'b010010001010110010: oled_data = 16'b1011001000101000;
				18'b010010001100110010: oled_data = 16'b1011001000001000;
				18'b010010001110110010: oled_data = 16'b1011001001101010;
				18'b010010010000110010: oled_data = 16'b1100011001011001;
				18'b010010010010110010: oled_data = 16'b1011111011111100;
				18'b010010010100110010: oled_data = 16'b1010011000111001;
				18'b010010010110110010: oled_data = 16'b1001010110110111;
				18'b010010011000110010: oled_data = 16'b1000110110110111;
				18'b010010011010110010: oled_data = 16'b1001110111111000;
				18'b010010011100110010: oled_data = 16'b1010111010011010;
				18'b010010011110110010: oled_data = 16'b1010101110101110;
				18'b010010100000110010: oled_data = 16'b1010000110100111;
				18'b010010100010110010: oled_data = 16'b1010000111000111;
				18'b010010100100110010: oled_data = 16'b1010000111000111;
				18'b010010100110110010: oled_data = 16'b1010000111000111;
				18'b010000011000110011: oled_data = 16'b1100110000110011;
				18'b010000011010110011: oled_data = 16'b1100110000010011;
				18'b010000011100110011: oled_data = 16'b1100110000110011;
				18'b010000011110110011: oled_data = 16'b1100110000110011;
				18'b010000100000110011: oled_data = 16'b1100110000110011;
				18'b010000100010110011: oled_data = 16'b1100110000110100;
				18'b010000100100110011: oled_data = 16'b1100001111110011;
				18'b010000100110110011: oled_data = 16'b1100110000010011;
				18'b010000101000110011: oled_data = 16'b1100001111110011;
				18'b010000101010110011: oled_data = 16'b1010001011001110;
				18'b010000101100110011: oled_data = 16'b1010001011101110;
				18'b010000101110110011: oled_data = 16'b1010001011101111;
				18'b010000110000110011: oled_data = 16'b1011001101010000;
				18'b010000110010110011: oled_data = 16'b1100110000010011;
				18'b010000110100110011: oled_data = 16'b1100110001010100;
				18'b010000110110110011: oled_data = 16'b1101010001010100;
				18'b010000111000110011: oled_data = 16'b1100110001010100;
				18'b010000111010110011: oled_data = 16'b1100110001010100;
				18'b010000111100110011: oled_data = 16'b1100110001010100;
				18'b010000111110110011: oled_data = 16'b1100110001010100;
				18'b010001000000110011: oled_data = 16'b1100110001010100;
				18'b010001000010110011: oled_data = 16'b1101010001010100;
				18'b010001000100110011: oled_data = 16'b1100010000010011;
				18'b010001000110110011: oled_data = 16'b1100010001010011;
				18'b010001001000110011: oled_data = 16'b1100010000110010;
				18'b010001001010110011: oled_data = 16'b1101010100010101;
				18'b010001001100110011: oled_data = 16'b1101111001111000;
				18'b010001001110110011: oled_data = 16'b1101111010111001;
				18'b010001010000110011: oled_data = 16'b1101111010111001;
				18'b010001010010110011: oled_data = 16'b1101111010111001;
				18'b010001010100110011: oled_data = 16'b1101111010111001;
				18'b010001010110110011: oled_data = 16'b1110011010111001;
				18'b010001011000110011: oled_data = 16'b1101111010111001;
				18'b010001011010110011: oled_data = 16'b1110011011011001;
				18'b010001011100110011: oled_data = 16'b1101011000110111;
				18'b010001011110110011: oled_data = 16'b1011110010110010;
				18'b010001100000110011: oled_data = 16'b1100010001010010;
				18'b010001100010110011: oled_data = 16'b1100010001010010;
				18'b010001100100110011: oled_data = 16'b1101010011010100;
				18'b010001100110110011: oled_data = 16'b1101010011010100;
				18'b010001101000110011: oled_data = 16'b1101010011010100;
				18'b010001101010110011: oled_data = 16'b1101010011010101;
				18'b010001101100110011: oled_data = 16'b1101010011010101;
				18'b010001101110110011: oled_data = 16'b1101010011010100;
				18'b010001110000110011: oled_data = 16'b1101010011010100;
				18'b010001110010110011: oled_data = 16'b1101110100110101;
				18'b010001110100110011: oled_data = 16'b1101111000111000;
				18'b010001110110110011: oled_data = 16'b1110011010111001;
				18'b010001111000110011: oled_data = 16'b1110011010111001;
				18'b010001111010110011: oled_data = 16'b1101111010011001;
				18'b010001111100110011: oled_data = 16'b1110011011011001;
				18'b010001111110110011: oled_data = 16'b1011001111001110;
				18'b010010000000110011: oled_data = 16'b1011001001001001;
				18'b010010000010110011: oled_data = 16'b1011101100001100;
				18'b010010000100110011: oled_data = 16'b1010101000001000;
				18'b010010000110110011: oled_data = 16'b1011001000001000;
				18'b010010001000110011: oled_data = 16'b1011001000001000;
				18'b010010001010110011: oled_data = 16'b1011001000001000;
				18'b010010001100110011: oled_data = 16'b1010101000001000;
				18'b010010001110110011: oled_data = 16'b1011001000001000;
				18'b010010010000110011: oled_data = 16'b1011110100010100;
				18'b010010010010110011: oled_data = 16'b1011011011111011;
				18'b010010010100110011: oled_data = 16'b1001010111010111;
				18'b010010010110110011: oled_data = 16'b1000110110010110;
				18'b010010011000110011: oled_data = 16'b1000110110010111;
				18'b010010011010110011: oled_data = 16'b1000110101110111;
				18'b010010011100110011: oled_data = 16'b1010010111010111;
				18'b010010011110110011: oled_data = 16'b1010001001101010;
				18'b010010100000110011: oled_data = 16'b1010000111000111;
				18'b010010100010110011: oled_data = 16'b1001100111000111;
				18'b010010100100110011: oled_data = 16'b1001100111000111;
				18'b010010100110110011: oled_data = 16'b1001100111000111;
				18'b010000011000110100: oled_data = 16'b1100101111110011;
				18'b010000011010110100: oled_data = 16'b1100101111110010;
				18'b010000011100110100: oled_data = 16'b1100110000010011;
				18'b010000011110110100: oled_data = 16'b1100110000010011;
				18'b010000100000110100: oled_data = 16'b1100110000010011;
				18'b010000100010110100: oled_data = 16'b1100101111110011;
				18'b010000100100110100: oled_data = 16'b1011101101110001;
				18'b010000100110110100: oled_data = 16'b1100110000010011;
				18'b010000101000110100: oled_data = 16'b1011001101010000;
				18'b010000101010110100: oled_data = 16'b1001101010101110;
				18'b010000101100110100: oled_data = 16'b1010001011101110;
				18'b010000101110110100: oled_data = 16'b1001101011001110;
				18'b010000110000110100: oled_data = 16'b1011101110010001;
				18'b010000110010110100: oled_data = 16'b1100010000010011;
				18'b010000110100110100: oled_data = 16'b1100110000110011;
				18'b010000110110110100: oled_data = 16'b1100110000110011;
				18'b010000111000110100: oled_data = 16'b1100110000110011;
				18'b010000111010110100: oled_data = 16'b1100110000110011;
				18'b010000111100110100: oled_data = 16'b1100110000110100;
				18'b010000111110110100: oled_data = 16'b1100110000110100;
				18'b010001000000110100: oled_data = 16'b1100110000110100;
				18'b010001000010110100: oled_data = 16'b1100110001010100;
				18'b010001000100110100: oled_data = 16'b1100010000010010;
				18'b010001000110110100: oled_data = 16'b1100110001110011;
				18'b010001001000110100: oled_data = 16'b1100010001010010;
				18'b010001001010110100: oled_data = 16'b1100110011110100;
				18'b010001001100110100: oled_data = 16'b1101011001011000;
				18'b010001001110110100: oled_data = 16'b1101111010011001;
				18'b010001010000110100: oled_data = 16'b1101111010111001;
				18'b010001010010110100: oled_data = 16'b1101111010111001;
				18'b010001010100110100: oled_data = 16'b1101111010111001;
				18'b010001010110110100: oled_data = 16'b1101111010111001;
				18'b010001011000110100: oled_data = 16'b1101111010111001;
				18'b010001011010110100: oled_data = 16'b1101111010111001;
				18'b010001011100110100: oled_data = 16'b1101111001111000;
				18'b010001011110110100: oled_data = 16'b1100110100110100;
				18'b010001100000110100: oled_data = 16'b1100110010110011;
				18'b010001100010110100: oled_data = 16'b1100110001110010;
				18'b010001100100110100: oled_data = 16'b1101010011010100;
				18'b010001100110110100: oled_data = 16'b1101010011010100;
				18'b010001101000110100: oled_data = 16'b1101010011010100;
				18'b010001101010110100: oled_data = 16'b1101010011010100;
				18'b010001101100110100: oled_data = 16'b1101010010110100;
				18'b010001101110110100: oled_data = 16'b1101010010110100;
				18'b010001110000110100: oled_data = 16'b1101010010110100;
				18'b010001110010110100: oled_data = 16'b1100010001110010;
				18'b010001110100110100: oled_data = 16'b1001110000010000;
				18'b010001110110110100: oled_data = 16'b1101011000010111;
				18'b010001111000110100: oled_data = 16'b1101011000010111;
				18'b010001111010110100: oled_data = 16'b1101010111110110;
				18'b010001111100110100: oled_data = 16'b1101111000110111;
				18'b010001111110110100: oled_data = 16'b1011001110001101;
				18'b010010000000110100: oled_data = 16'b1011001000101000;
				18'b010010000010110100: oled_data = 16'b1011001011001011;
				18'b010010000100110100: oled_data = 16'b1010101000001000;
				18'b010010000110110100: oled_data = 16'b1010101000001000;
				18'b010010001000110100: oled_data = 16'b1010101000001000;
				18'b010010001010110100: oled_data = 16'b1010101000001000;
				18'b010010001100110100: oled_data = 16'b1010101000001000;
				18'b010010001110110100: oled_data = 16'b1010101000001000;
				18'b010010010000110100: oled_data = 16'b1001101001001010;
				18'b010010010010110100: oled_data = 16'b1011111000011000;
				18'b010010010100110100: oled_data = 16'b1001111000111000;
				18'b010010010110110100: oled_data = 16'b1000110110010110;
				18'b010010011000110100: oled_data = 16'b1000110110010111;
				18'b010010011010110100: oled_data = 16'b1001010110110111;
				18'b010010011100110100: oled_data = 16'b1010001110101111;
				18'b010010011110110100: oled_data = 16'b1001100110100111;
				18'b010010100000110100: oled_data = 16'b1010000111000111;
				18'b010010100010110100: oled_data = 16'b1001100111000111;
				18'b010010100100110100: oled_data = 16'b1001100110100111;
				18'b010010100110110100: oled_data = 16'b1001100110100111;
				18'b010000011000110101: oled_data = 16'b1100101111010010;
				18'b010000011010110101: oled_data = 16'b1100101111010010;
				18'b010000011100110101: oled_data = 16'b1100001111010010;
				18'b010000011110110101: oled_data = 16'b1100001111010010;
				18'b010000100000110101: oled_data = 16'b1100001111110010;
				18'b010000100010110101: oled_data = 16'b1011001101110000;
				18'b010000100100110101: oled_data = 16'b1011001101110000;
				18'b010000100110110101: oled_data = 16'b1100001111110010;
				18'b010000101000110101: oled_data = 16'b1010001011001110;
				18'b010000101010110101: oled_data = 16'b1001101010101110;
				18'b010000101100110101: oled_data = 16'b1001101011001110;
				18'b010000101110110101: oled_data = 16'b1001101010101101;
				18'b010000110000110101: oled_data = 16'b1011101110110001;
				18'b010000110010110101: oled_data = 16'b1100001111010010;
				18'b010000110100110101: oled_data = 16'b1100101111110011;
				18'b010000110110110101: oled_data = 16'b1100101111110011;
				18'b010000111000110101: oled_data = 16'b1100101111110011;
				18'b010000111010110101: oled_data = 16'b1100110000010011;
				18'b010000111100110101: oled_data = 16'b1100110000010011;
				18'b010000111110110101: oled_data = 16'b1100110000010011;
				18'b010001000000110101: oled_data = 16'b1100110000010011;
				18'b010001000010110101: oled_data = 16'b1100110000010011;
				18'b010001000100110101: oled_data = 16'b1100001111110010;
				18'b010001000110110101: oled_data = 16'b1011110000010010;
				18'b010001001000110101: oled_data = 16'b1100010001010010;
				18'b010001001010110101: oled_data = 16'b1100110100110101;
				18'b010001001100110101: oled_data = 16'b1101011001111000;
				18'b010001001110110101: oled_data = 16'b1101111010011000;
				18'b010001010000110101: oled_data = 16'b1101111010011000;
				18'b010001010010110101: oled_data = 16'b1101111010011000;
				18'b010001010100110101: oled_data = 16'b1101111010011000;
				18'b010001010110110101: oled_data = 16'b1101111010011001;
				18'b010001011000110101: oled_data = 16'b1101111010011000;
				18'b010001011010110101: oled_data = 16'b1101111010011001;
				18'b010001011100110101: oled_data = 16'b1101111001111000;
				18'b010001011110110101: oled_data = 16'b1100110101010101;
				18'b010001100000110101: oled_data = 16'b1100110001110010;
				18'b010001100010110101: oled_data = 16'b1100010000110001;
				18'b010001100100110101: oled_data = 16'b1101010010110011;
				18'b010001100110110101: oled_data = 16'b1101010010110011;
				18'b010001101000110101: oled_data = 16'b1101010010110011;
				18'b010001101010110101: oled_data = 16'b1101010010110011;
				18'b010001101100110101: oled_data = 16'b1101010010010100;
				18'b010001101110110101: oled_data = 16'b1101010010110100;
				18'b010001110000110101: oled_data = 16'b1101010010110100;
				18'b010001110010110101: oled_data = 16'b1010101110101111;
				18'b010001110100110101: oled_data = 16'b0010100010100010;
				18'b010001110110110101: oled_data = 16'b0110101011101011;
				18'b010001111000110101: oled_data = 16'b1010110010110010;
				18'b010001111010110101: oled_data = 16'b1011010011010010;
				18'b010001111100110101: oled_data = 16'b1011110011010011;
				18'b010001111110110101: oled_data = 16'b1010001010101011;
				18'b010010000000110101: oled_data = 16'b1010100111101000;
				18'b010010000010110101: oled_data = 16'b1011001010101010;
				18'b010010000100110101: oled_data = 16'b1010101000001000;
				18'b010010000110110101: oled_data = 16'b1010101000001000;
				18'b010010001000110101: oled_data = 16'b1010101000001000;
				18'b010010001010110101: oled_data = 16'b1010101000001000;
				18'b010010001100110101: oled_data = 16'b1010100111101000;
				18'b010010001110110101: oled_data = 16'b1010000111101000;
				18'b010010010000110101: oled_data = 16'b1000100101000110;
				18'b010010010010110101: oled_data = 16'b1010101011001100;
				18'b010010010100110101: oled_data = 16'b1011010011010011;
				18'b010010010110110101: oled_data = 16'b1010010011010100;
				18'b010010011000110101: oled_data = 16'b1010010001010010;
				18'b010010011010110101: oled_data = 16'b1010001101001110;
				18'b010010011100110101: oled_data = 16'b1001100111000111;
				18'b010010011110110101: oled_data = 16'b1010000111000111;
				18'b010010100000110101: oled_data = 16'b1001100111000111;
				18'b010010100010110101: oled_data = 16'b1001100110100111;
				18'b010010100100110101: oled_data = 16'b1001100110100111;
				18'b010010100110110101: oled_data = 16'b1001100110100111;
				18'b010000011000110110: oled_data = 16'b1100001111010010;
				18'b010000011010110110: oled_data = 16'b1100001110110010;
				18'b010000011100110110: oled_data = 16'b1100001110110010;
				18'b010000011110110110: oled_data = 16'b1100001110110010;
				18'b010000100000110110: oled_data = 16'b1011101110010001;
				18'b010000100010110110: oled_data = 16'b1010001011001110;
				18'b010000100100110110: oled_data = 16'b1100001111010010;
				18'b010000100110110110: oled_data = 16'b1011001101010000;
				18'b010000101000110110: oled_data = 16'b1001001001101101;
				18'b010000101010110110: oled_data = 16'b1001101010001101;
				18'b010000101100110110: oled_data = 16'b1001101010001101;
				18'b010000101110110110: oled_data = 16'b1001101011001110;
				18'b010000110000110110: oled_data = 16'b1100001111010010;
				18'b010000110010110110: oled_data = 16'b1100001111010010;
				18'b010000110100110110: oled_data = 16'b1100001111010010;
				18'b010000110110110110: oled_data = 16'b1100101111010010;
				18'b010000111000110110: oled_data = 16'b1100101111110010;
				18'b010000111010110110: oled_data = 16'b1100101111110010;
				18'b010000111100110110: oled_data = 16'b1100101111110011;
				18'b010000111110110110: oled_data = 16'b1100101111110011;
				18'b010001000000110110: oled_data = 16'b1100101111110011;
				18'b010001000010110110: oled_data = 16'b1100001111110010;
				18'b010001000100110110: oled_data = 16'b1100010000010010;
				18'b010001000110110110: oled_data = 16'b1100010000010010;
				18'b010001001000110110: oled_data = 16'b1100010001010010;
				18'b010001001010110110: oled_data = 16'b1100110101010101;
				18'b010001001100110110: oled_data = 16'b1101011001011000;
				18'b010001001110110110: oled_data = 16'b1101011001111000;
				18'b010001010000110110: oled_data = 16'b1101011001111000;
				18'b010001010010110110: oled_data = 16'b1101011001111000;
				18'b010001010100110110: oled_data = 16'b1101011001111000;
				18'b010001010110110110: oled_data = 16'b1101111001111000;
				18'b010001011000110110: oled_data = 16'b1101011001111000;
				18'b010001011010110110: oled_data = 16'b1101011001011000;
				18'b010001011100110110: oled_data = 16'b1101011000110111;
				18'b010001011110110110: oled_data = 16'b1100010100110100;
				18'b010001100000110110: oled_data = 16'b1100010001010010;
				18'b010001100010110110: oled_data = 16'b1100010000110010;
				18'b010001100100110110: oled_data = 16'b1100110010010011;
				18'b010001100110110110: oled_data = 16'b1100110010010011;
				18'b010001101000110110: oled_data = 16'b1100110010010011;
				18'b010001101010110110: oled_data = 16'b1100110010010011;
				18'b010001101100110110: oled_data = 16'b1100110010010011;
				18'b010001101110110110: oled_data = 16'b1100110010010011;
				18'b010001110000110110: oled_data = 16'b1101010010010100;
				18'b010001110010110110: oled_data = 16'b0110101000001001;
				18'b010001110100110110: oled_data = 16'b0010000001100001;
				18'b010001110110110110: oled_data = 16'b0010100010100010;
				18'b010001111000110110: oled_data = 16'b0100100110000101;
				18'b010001111010110110: oled_data = 16'b1000001011001011;
				18'b010001111100110110: oled_data = 16'b1010001110101111;
				18'b010001111110110110: oled_data = 16'b1001101010001010;
				18'b010010000000110110: oled_data = 16'b1010100111101000;
				18'b010010000010110110: oled_data = 16'b1010101001101001;
				18'b010010000100110110: oled_data = 16'b1010100111101000;
				18'b010010000110110110: oled_data = 16'b1010100111101000;
				18'b010010001000110110: oled_data = 16'b1010100111101000;
				18'b010010001010110110: oled_data = 16'b1010000111101000;
				18'b010010001100110110: oled_data = 16'b1010100111100111;
				18'b010010001110110110: oled_data = 16'b1001100111000111;
				18'b010010010000110110: oled_data = 16'b1000100110000110;
				18'b010010010010110110: oled_data = 16'b1010000111000111;
				18'b010010010100110110: oled_data = 16'b1010000111000111;
				18'b010010010110110110: oled_data = 16'b1010000111101000;
				18'b010010011000110110: oled_data = 16'b1001100110100111;
				18'b010010011010110110: oled_data = 16'b1010000110100111;
				18'b010010011100110110: oled_data = 16'b1010000111000111;
				18'b010010011110110110: oled_data = 16'b1001100110100111;
				18'b010010100000110110: oled_data = 16'b1001100110100111;
				18'b010010100010110110: oled_data = 16'b1001100110100110;
				18'b010010100100110110: oled_data = 16'b1001000110000110;
				18'b010010100110110110: oled_data = 16'b1001000110000110;
				18'b010000011000110111: oled_data = 16'b1100001110110001;
				18'b010000011010110111: oled_data = 16'b1100001110110001;
				18'b010000011100110111: oled_data = 16'b1100001110110001;
				18'b010000011110110111: oled_data = 16'b1100001110110001;
				18'b010000100000110111: oled_data = 16'b1010001011001110;
				18'b010000100010110111: oled_data = 16'b1001101010101101;
				18'b010000100100110111: oled_data = 16'b1100001111010010;
				18'b010000100110110111: oled_data = 16'b1010001011001110;
				18'b010000101000110111: oled_data = 16'b1001001001101101;
				18'b010000101010110111: oled_data = 16'b1001001010001101;
				18'b010000101100110111: oled_data = 16'b1001001010001101;
				18'b010000101110110111: oled_data = 16'b1010001011001110;
				18'b010000110000110111: oled_data = 16'b1100001111010001;
				18'b010000110010110111: oled_data = 16'b1100001110110001;
				18'b010000110100110111: oled_data = 16'b1011101110110001;
				18'b010000110110110111: oled_data = 16'b1100001111010010;
				18'b010000111000110111: oled_data = 16'b1100001111010010;
				18'b010000111010110111: oled_data = 16'b1100001111010010;
				18'b010000111100110111: oled_data = 16'b1100001111010010;
				18'b010000111110110111: oled_data = 16'b1100001111010010;
				18'b010001000000110111: oled_data = 16'b1100001111010010;
				18'b010001000010110111: oled_data = 16'b1100001111010010;
				18'b010001000100110111: oled_data = 16'b1100110000010011;
				18'b010001000110110111: oled_data = 16'b1100110000110011;
				18'b010001001000110111: oled_data = 16'b1100110000110010;
				18'b010001001010110111: oled_data = 16'b1100110101110101;
				18'b010001001100110111: oled_data = 16'b1101011001010111;
				18'b010001001110110111: oled_data = 16'b1101011001010111;
				18'b010001010000110111: oled_data = 16'b1101011001010111;
				18'b010001010010110111: oled_data = 16'b1101011001010111;
				18'b010001010100110111: oled_data = 16'b1101011001010111;
				18'b010001010110110111: oled_data = 16'b1101011001010111;
				18'b010001011000110111: oled_data = 16'b1101011000110111;
				18'b010001011010110111: oled_data = 16'b1101011001010111;
				18'b010001011100110111: oled_data = 16'b1101010111110110;
				18'b010001011110110111: oled_data = 16'b1100010011110011;
				18'b010001100000110111: oled_data = 16'b1100010001010010;
				18'b010001100010110111: oled_data = 16'b1100010000110010;
				18'b010001100100110111: oled_data = 16'b1100110001110010;
				18'b010001100110110111: oled_data = 16'b1100110001110010;
				18'b010001101000110111: oled_data = 16'b1100110001110010;
				18'b010001101010110111: oled_data = 16'b1100110001110010;
				18'b010001101100110111: oled_data = 16'b1100110001110010;
				18'b010001101110110111: oled_data = 16'b1100110001110011;
				18'b010001110000110111: oled_data = 16'b1011110000010001;
				18'b010001110010110111: oled_data = 16'b0011100010100011;
				18'b010001110100110111: oled_data = 16'b0011100011100010;
				18'b010001110110110111: oled_data = 16'b0101000110000100;
				18'b010001111000110111: oled_data = 16'b0110101001000111;
				18'b010001111010110111: oled_data = 16'b0111101001000111;
				18'b010001111100110111: oled_data = 16'b1000001001100111;
				18'b010001111110110111: oled_data = 16'b1000101000000111;
				18'b010010000000110111: oled_data = 16'b1010100111101000;
				18'b010010000010110111: oled_data = 16'b1010001000101000;
				18'b010010000100110111: oled_data = 16'b1010100111101000;
				18'b010010000110110111: oled_data = 16'b1010100111100111;
				18'b010010001000110111: oled_data = 16'b1010000111100111;
				18'b010010001010110111: oled_data = 16'b1010000111100111;
				18'b010010001100110111: oled_data = 16'b1010000111000111;
				18'b010010001110110111: oled_data = 16'b1001100110100111;
				18'b010010010000110111: oled_data = 16'b1000100110000111;
				18'b010010010010110111: oled_data = 16'b1010000111001000;
				18'b010010010100110111: oled_data = 16'b1010000111000111;
				18'b010010010110110111: oled_data = 16'b1001100110100111;
				18'b010010011000110111: oled_data = 16'b1001000110100110;
				18'b010010011010110111: oled_data = 16'b1001100110100111;
				18'b010010011100110111: oled_data = 16'b1001100110100111;
				18'b010010011110110111: oled_data = 16'b1001100110100110;
				18'b010010100000110111: oled_data = 16'b1001100110000110;
				18'b010010100010110111: oled_data = 16'b1001000110000110;
				18'b010010100100110111: oled_data = 16'b1001000110000110;
				18'b010010100110110111: oled_data = 16'b1001000110000110;
				18'b010100011000001000: oled_data = 16'b1001101111101011;
				18'b010100011010001000: oled_data = 16'b1010010000001011;
				18'b010100011100001000: oled_data = 16'b1010010000101011;
				18'b010100011110001000: oled_data = 16'b1010110001001100;
				18'b010100100000001000: oled_data = 16'b1010110000001011;
				18'b010100100010001000: oled_data = 16'b1101110111110110;
				18'b010100100100001000: oled_data = 16'b1111011010011100;
				18'b010100100110001000: oled_data = 16'b1110010100010110;
				18'b010100101000001000: oled_data = 16'b1101110010110101;
				18'b010100101010001000: oled_data = 16'b1101110011010101;
				18'b010100101100001000: oled_data = 16'b1101110011010101;
				18'b010100101110001000: oled_data = 16'b1101110011010101;
				18'b010100110000001000: oled_data = 16'b1101110011010101;
				18'b010100110010001000: oled_data = 16'b1101110011010101;
				18'b010100110100001000: oled_data = 16'b1101110011010101;
				18'b010100110110001000: oled_data = 16'b1101110011010101;
				18'b010100111000001000: oled_data = 16'b1101110011010101;
				18'b010100111010001000: oled_data = 16'b1101110011010101;
				18'b010100111100001000: oled_data = 16'b1101110011010101;
				18'b010100111110001000: oled_data = 16'b1101110011010101;
				18'b010101000000001000: oled_data = 16'b1101110011010101;
				18'b010101000010001000: oled_data = 16'b1101110011010101;
				18'b010101000100001000: oled_data = 16'b1101110011010101;
				18'b010101000110001000: oled_data = 16'b1101110011010101;
				18'b010101001000001000: oled_data = 16'b1101110011010101;
				18'b010101001010001000: oled_data = 16'b1101110011010101;
				18'b010101001100001000: oled_data = 16'b1101110011010101;
				18'b010101001110001000: oled_data = 16'b1101110011010101;
				18'b010101010000001000: oled_data = 16'b1101110011010101;
				18'b010101010010001000: oled_data = 16'b1101110011010101;
				18'b010101010100001000: oled_data = 16'b1101110011010101;
				18'b010101010110001000: oled_data = 16'b1101110011010101;
				18'b010101011000001000: oled_data = 16'b1101110011010101;
				18'b010101011010001000: oled_data = 16'b1101110011010101;
				18'b010101011100001000: oled_data = 16'b1101110011010101;
				18'b010101011110001000: oled_data = 16'b1101110011010101;
				18'b010101100000001000: oled_data = 16'b1101110011010101;
				18'b010101100010001000: oled_data = 16'b1101110011010101;
				18'b010101100100001000: oled_data = 16'b1101110011010101;
				18'b010101100110001000: oled_data = 16'b1101110011010101;
				18'b010101101000001000: oled_data = 16'b1101110011010101;
				18'b010101101010001000: oled_data = 16'b1101110011010101;
				18'b010101101100001000: oled_data = 16'b1101110011010101;
				18'b010101101110001000: oled_data = 16'b1110010011010110;
				18'b010101110000001000: oled_data = 16'b1101110010110101;
				18'b010101110010001000: oled_data = 16'b1101010010010100;
				18'b010101110100001000: oled_data = 16'b1101110011010110;
				18'b010101110110001000: oled_data = 16'b1101110011010101;
				18'b010101111000001000: oled_data = 16'b1101110011010110;
				18'b010101111010001000: oled_data = 16'b1101010010010100;
				18'b010101111100001000: oled_data = 16'b1101010010010100;
				18'b010101111110001000: oled_data = 16'b1101110011010101;
				18'b010110000000001000: oled_data = 16'b1101110011010101;
				18'b010110000010001000: oled_data = 16'b1101010010110101;
				18'b010110000100001000: oled_data = 16'b1110111000111010;
				18'b010110000110001000: oled_data = 16'b1101111000111001;
				18'b010110001000001000: oled_data = 16'b0101101001000111;
				18'b010110001010001000: oled_data = 16'b0101101001000101;
				18'b010110001100001000: oled_data = 16'b0111001011000110;
				18'b010110001110001000: oled_data = 16'b0111101011100111;
				18'b010110010000001000: oled_data = 16'b0111101100000111;
				18'b010110010010001000: oled_data = 16'b0111101100000111;
				18'b010110010100001000: oled_data = 16'b0111001100000111;
				18'b010110010110001000: oled_data = 16'b0111001011101000;
				18'b010110011000001000: oled_data = 16'b0110101011101000;
				18'b010110011010001000: oled_data = 16'b0110001011001000;
				18'b010110011100001000: oled_data = 16'b0110001010101000;
				18'b010110011110001000: oled_data = 16'b0101101010001000;
				18'b010110100000001000: oled_data = 16'b0101101010001000;
				18'b010110100010001000: oled_data = 16'b0101001001101000;
				18'b010110100100001000: oled_data = 16'b0101001001001000;
				18'b010110100110001000: oled_data = 16'b0101001001101000;
				18'b010100011000001001: oled_data = 16'b1011010001101011;
				18'b010100011010001001: oled_data = 16'b1011010001101011;
				18'b010100011100001001: oled_data = 16'b1011010001001011;
				18'b010100011110001001: oled_data = 16'b1010110000101011;
				18'b010100100000001001: oled_data = 16'b1011110010101111;
				18'b010100100010001001: oled_data = 16'b1111011010111011;
				18'b010100100100001001: oled_data = 16'b1110010111011000;
				18'b010100100110001001: oled_data = 16'b1101110011010101;
				18'b010100101000001001: oled_data = 16'b1101110011010101;
				18'b010100101010001001: oled_data = 16'b1101110011010101;
				18'b010100101100001001: oled_data = 16'b1101110011010101;
				18'b010100101110001001: oled_data = 16'b1101110011010101;
				18'b010100110000001001: oled_data = 16'b1101110011010101;
				18'b010100110010001001: oled_data = 16'b1101110011010101;
				18'b010100110100001001: oled_data = 16'b1101110011010101;
				18'b010100110110001001: oled_data = 16'b1101110011010101;
				18'b010100111000001001: oled_data = 16'b1101110011010101;
				18'b010100111010001001: oled_data = 16'b1101110011010101;
				18'b010100111100001001: oled_data = 16'b1101110011010101;
				18'b010100111110001001: oled_data = 16'b1101110011010101;
				18'b010101000000001001: oled_data = 16'b1101110011010101;
				18'b010101000010001001: oled_data = 16'b1101110011010101;
				18'b010101000100001001: oled_data = 16'b1101110011010101;
				18'b010101000110001001: oled_data = 16'b1101110011010101;
				18'b010101001000001001: oled_data = 16'b1101110011010101;
				18'b010101001010001001: oled_data = 16'b1101110011010101;
				18'b010101001100001001: oled_data = 16'b1101110011010101;
				18'b010101001110001001: oled_data = 16'b1101110011010101;
				18'b010101010000001001: oled_data = 16'b1101110011010101;
				18'b010101010010001001: oled_data = 16'b1101110011010101;
				18'b010101010100001001: oled_data = 16'b1101110011010101;
				18'b010101010110001001: oled_data = 16'b1101110011010110;
				18'b010101011000001001: oled_data = 16'b1101110010010101;
				18'b010101011010001001: oled_data = 16'b1101110010110101;
				18'b010101011100001001: oled_data = 16'b1101110011010101;
				18'b010101011110001001: oled_data = 16'b1101110011010101;
				18'b010101100000001001: oled_data = 16'b1101110011010101;
				18'b010101100010001001: oled_data = 16'b1101110011010101;
				18'b010101100100001001: oled_data = 16'b1101110011010101;
				18'b010101100110001001: oled_data = 16'b1101110011010101;
				18'b010101101000001001: oled_data = 16'b1101110011010101;
				18'b010101101010001001: oled_data = 16'b1101010001110100;
				18'b010101101100001001: oled_data = 16'b1101110011010101;
				18'b010101101110001001: oled_data = 16'b1101110011010110;
				18'b010101110000001001: oled_data = 16'b1101110011010110;
				18'b010101110010001001: oled_data = 16'b1101010010010100;
				18'b010101110100001001: oled_data = 16'b1101110011010101;
				18'b010101110110001001: oled_data = 16'b1101110011010101;
				18'b010101111000001001: oled_data = 16'b1110010011010110;
				18'b010101111010001001: oled_data = 16'b1101110011010101;
				18'b010101111100001001: oled_data = 16'b1101010010010100;
				18'b010101111110001001: oled_data = 16'b1101110011010101;
				18'b010110000000001001: oled_data = 16'b1101110011010101;
				18'b010110000010001001: oled_data = 16'b1101010010110101;
				18'b010110000100001001: oled_data = 16'b1101010101010110;
				18'b010110000110001001: oled_data = 16'b1111011100011101;
				18'b010110001000001001: oled_data = 16'b1000101111001101;
				18'b010110001010001001: oled_data = 16'b0101101000100101;
				18'b010110001100001001: oled_data = 16'b0111001011000110;
				18'b010110001110001001: oled_data = 16'b0111101011100111;
				18'b010110010000001001: oled_data = 16'b0111101100000111;
				18'b010110010010001001: oled_data = 16'b1000001100100111;
				18'b010110010100001001: oled_data = 16'b1000001100100111;
				18'b010110010110001001: oled_data = 16'b1000101101001000;
				18'b010110011000001001: oled_data = 16'b1000101101101000;
				18'b010110011010001001: oled_data = 16'b1000101101101000;
				18'b010110011100001001: oled_data = 16'b1000101101101000;
				18'b010110011110001001: oled_data = 16'b1000101110001001;
				18'b010110100000001001: oled_data = 16'b1000101110101010;
				18'b010110100010001001: oled_data = 16'b0101101010101000;
				18'b010110100100001001: oled_data = 16'b0011101000000111;
				18'b010110100110001001: oled_data = 16'b0100001000101000;
				18'b010100011000001010: oled_data = 16'b1011010001101100;
				18'b010100011010001010: oled_data = 16'b1011010001101011;
				18'b010100011100001010: oled_data = 16'b1011010001001011;
				18'b010100011110001010: oled_data = 16'b1010110000101011;
				18'b010100100000001010: oled_data = 16'b1101010111010101;
				18'b010100100010001010: oled_data = 16'b1111011001111011;
				18'b010100100100001010: oled_data = 16'b1110010100010110;
				18'b010100100110001010: oled_data = 16'b1101110011010101;
				18'b010100101000001010: oled_data = 16'b1101110011010101;
				18'b010100101010001010: oled_data = 16'b1101110011010101;
				18'b010100101100001010: oled_data = 16'b1101110011010101;
				18'b010100101110001010: oled_data = 16'b1101110011010101;
				18'b010100110000001010: oled_data = 16'b1101110011010101;
				18'b010100110010001010: oled_data = 16'b1101110011010101;
				18'b010100110100001010: oled_data = 16'b1101110011010101;
				18'b010100110110001010: oled_data = 16'b1101110010110101;
				18'b010100111000001010: oled_data = 16'b1101110011010101;
				18'b010100111010001010: oled_data = 16'b1101110011010101;
				18'b010100111100001010: oled_data = 16'b1101110011010101;
				18'b010100111110001010: oled_data = 16'b1101110011010101;
				18'b010101000000001010: oled_data = 16'b1101110011010101;
				18'b010101000010001010: oled_data = 16'b1101110011010101;
				18'b010101000100001010: oled_data = 16'b1101110011010101;
				18'b010101000110001010: oled_data = 16'b1101110011010101;
				18'b010101001000001010: oled_data = 16'b1101110011010101;
				18'b010101001010001010: oled_data = 16'b1101110011010101;
				18'b010101001100001010: oled_data = 16'b1101110011010101;
				18'b010101001110001010: oled_data = 16'b1101110011010101;
				18'b010101010000001010: oled_data = 16'b1101110011010101;
				18'b010101010010001010: oled_data = 16'b1101110011010101;
				18'b010101010100001010: oled_data = 16'b1101110011010101;
				18'b010101010110001010: oled_data = 16'b1101110011010110;
				18'b010101011000001010: oled_data = 16'b1101010010010100;
				18'b010101011010001010: oled_data = 16'b1101110010110101;
				18'b010101011100001010: oled_data = 16'b1101110011010101;
				18'b010101011110001010: oled_data = 16'b1101110011010101;
				18'b010101100000001010: oled_data = 16'b1101110011010101;
				18'b010101100010001010: oled_data = 16'b1101110011010101;
				18'b010101100100001010: oled_data = 16'b1101110011010101;
				18'b010101100110001010: oled_data = 16'b1101110011010101;
				18'b010101101000001010: oled_data = 16'b1101110011010110;
				18'b010101101010001010: oled_data = 16'b1101110010010101;
				18'b010101101100001010: oled_data = 16'b1101110010110101;
				18'b010101101110001010: oled_data = 16'b1101110011010110;
				18'b010101110000001010: oled_data = 16'b1101110011010110;
				18'b010101110010001010: oled_data = 16'b1101010010010101;
				18'b010101110100001010: oled_data = 16'b1101110010010101;
				18'b010101110110001010: oled_data = 16'b1110010011010110;
				18'b010101111000001010: oled_data = 16'b1110010011010110;
				18'b010101111010001010: oled_data = 16'b1101110011010110;
				18'b010101111100001010: oled_data = 16'b1101010010010100;
				18'b010101111110001010: oled_data = 16'b1101110011010101;
				18'b010110000000001010: oled_data = 16'b1101110011010101;
				18'b010110000010001010: oled_data = 16'b1101110010110101;
				18'b010110000100001010: oled_data = 16'b1101010011110110;
				18'b010110000110001010: oled_data = 16'b1111011011111100;
				18'b010110001000001010: oled_data = 16'b1100010101110110;
				18'b010110001010001010: oled_data = 16'b0011100101100101;
				18'b010110001100001010: oled_data = 16'b0100000111000110;
				18'b010110001110001010: oled_data = 16'b0101001000000110;
				18'b010110010000001010: oled_data = 16'b0101101001000110;
				18'b010110010010001010: oled_data = 16'b0110101010100111;
				18'b010110010100001010: oled_data = 16'b0111101011101000;
				18'b010110010110001010: oled_data = 16'b0111101100001000;
				18'b010110011000001010: oled_data = 16'b1000101101001000;
				18'b010110011010001010: oled_data = 16'b1000101101101000;
				18'b010110011100001010: oled_data = 16'b1000101110001000;
				18'b010110011110001010: oled_data = 16'b1000101110001000;
				18'b010110100000001010: oled_data = 16'b1000101110001001;
				18'b010110100010001010: oled_data = 16'b0111001011101001;
				18'b010110100100001010: oled_data = 16'b1001001101001101;
				18'b010110100110001010: oled_data = 16'b1011110000010001;
				18'b010100011000001011: oled_data = 16'b1001001111001010;
				18'b010100011010001011: oled_data = 16'b1000101110001001;
				18'b010100011100001011: oled_data = 16'b0111101100001001;
				18'b010100011110001011: oled_data = 16'b1000101110101100;
				18'b010100100000001011: oled_data = 16'b1110111001111010;
				18'b010100100010001011: oled_data = 16'b1110010110111001;
				18'b010100100100001011: oled_data = 16'b1101110011010101;
				18'b010100100110001011: oled_data = 16'b1101110011010101;
				18'b010100101000001011: oled_data = 16'b1101110011010101;
				18'b010100101010001011: oled_data = 16'b1101110011010101;
				18'b010100101100001011: oled_data = 16'b1101110011010101;
				18'b010100101110001011: oled_data = 16'b1101110011010101;
				18'b010100110000001011: oled_data = 16'b1101110011010101;
				18'b010100110010001011: oled_data = 16'b1101110011010101;
				18'b010100110100001011: oled_data = 16'b1101110010110101;
				18'b010100110110001011: oled_data = 16'b1101010010010100;
				18'b010100111000001011: oled_data = 16'b1101110011010110;
				18'b010100111010001011: oled_data = 16'b1101110011010101;
				18'b010100111100001011: oled_data = 16'b1101110011010101;
				18'b010100111110001011: oled_data = 16'b1101110011010101;
				18'b010101000000001011: oled_data = 16'b1101110011010101;
				18'b010101000010001011: oled_data = 16'b1101110011010101;
				18'b010101000100001011: oled_data = 16'b1101110011010101;
				18'b010101000110001011: oled_data = 16'b1101110011010101;
				18'b010101001000001011: oled_data = 16'b1101110011010101;
				18'b010101001010001011: oled_data = 16'b1101110011010101;
				18'b010101001100001011: oled_data = 16'b1101110011010101;
				18'b010101001110001011: oled_data = 16'b1101110011010101;
				18'b010101010000001011: oled_data = 16'b1101110011010101;
				18'b010101010010001011: oled_data = 16'b1101110011010101;
				18'b010101010100001011: oled_data = 16'b1101110011010101;
				18'b010101010110001011: oled_data = 16'b1101110011010101;
				18'b010101011000001011: oled_data = 16'b1101010010010100;
				18'b010101011010001011: oled_data = 16'b1101110011010101;
				18'b010101011100001011: oled_data = 16'b1101110011010101;
				18'b010101011110001011: oled_data = 16'b1101110011010101;
				18'b010101100000001011: oled_data = 16'b1101110011010101;
				18'b010101100010001011: oled_data = 16'b1101110011010101;
				18'b010101100100001011: oled_data = 16'b1101110011010101;
				18'b010101100110001011: oled_data = 16'b1110010011010110;
				18'b010101101000001011: oled_data = 16'b1110010011110110;
				18'b010101101010001011: oled_data = 16'b1101110010110101;
				18'b010101101100001011: oled_data = 16'b1101010010010100;
				18'b010101101110001011: oled_data = 16'b1101110011010110;
				18'b010101110000001011: oled_data = 16'b1101110011010101;
				18'b010101110010001011: oled_data = 16'b1101110010110101;
				18'b010101110100001011: oled_data = 16'b1101010001110100;
				18'b010101110110001011: oled_data = 16'b1101110011010110;
				18'b010101111000001011: oled_data = 16'b1101110011010101;
				18'b010101111010001011: oled_data = 16'b1110010011010110;
				18'b010101111100001011: oled_data = 16'b1101010010010100;
				18'b010101111110001011: oled_data = 16'b1101110010110101;
				18'b010110000000001011: oled_data = 16'b1101110011010101;
				18'b010110000010001011: oled_data = 16'b1101110011010101;
				18'b010110000100001011: oled_data = 16'b1101010011010101;
				18'b010110000110001011: oled_data = 16'b1110111000111010;
				18'b010110001000001011: oled_data = 16'b1110111010111011;
				18'b010110001010001011: oled_data = 16'b0100000111000111;
				18'b010110001100001011: oled_data = 16'b0010000100100101;
				18'b010110001110001011: oled_data = 16'b0010000101000101;
				18'b010110010000001011: oled_data = 16'b0010000101100110;
				18'b010110010010001011: oled_data = 16'b0010100110000110;
				18'b010110010100001011: oled_data = 16'b0011100111000110;
				18'b010110010110001011: oled_data = 16'b0100001000000111;
				18'b010110011000001011: oled_data = 16'b0101001000100111;
				18'b010110011010001011: oled_data = 16'b0101101001100111;
				18'b010110011100001011: oled_data = 16'b0111001011001000;
				18'b010110011110001011: oled_data = 16'b1010001110001100;
				18'b010110100000001011: oled_data = 16'b1100010001010000;
				18'b010110100010001011: oled_data = 16'b1101110010110010;
				18'b010110100100001011: oled_data = 16'b1101110001010001;
				18'b010110100110001011: oled_data = 16'b1100101101101110;
				18'b010100011000001100: oled_data = 16'b0101101011001000;
				18'b010100011010001100: oled_data = 16'b0110001010101000;
				18'b010100011100001100: oled_data = 16'b0111001010101000;
				18'b010100011110001100: oled_data = 16'b1011010011010010;
				18'b010100100000001100: oled_data = 16'b1111011010111011;
				18'b010100100010001100: oled_data = 16'b1110010100010110;
				18'b010100100100001100: oled_data = 16'b1101110011010110;
				18'b010100100110001100: oled_data = 16'b1101110011010110;
				18'b010100101000001100: oled_data = 16'b1101110011010101;
				18'b010100101010001100: oled_data = 16'b1101110011010101;
				18'b010100101100001100: oled_data = 16'b1101110011010101;
				18'b010100101110001100: oled_data = 16'b1101110011010101;
				18'b010100110000001100: oled_data = 16'b1101110011010101;
				18'b010100110010001100: oled_data = 16'b1101110011010101;
				18'b010100110100001100: oled_data = 16'b1101010010010100;
				18'b010100110110001100: oled_data = 16'b1101110011010101;
				18'b010100111000001100: oled_data = 16'b1101110011010101;
				18'b010100111010001100: oled_data = 16'b1101110011010101;
				18'b010100111100001100: oled_data = 16'b1101110011010110;
				18'b010100111110001100: oled_data = 16'b1101110011010101;
				18'b010101000000001100: oled_data = 16'b1101110011010101;
				18'b010101000010001100: oled_data = 16'b1101110011010101;
				18'b010101000100001100: oled_data = 16'b1101110011010101;
				18'b010101000110001100: oled_data = 16'b1101110011010101;
				18'b010101001000001100: oled_data = 16'b1101110011010101;
				18'b010101001010001100: oled_data = 16'b1101110011010101;
				18'b010101001100001100: oled_data = 16'b1101110011010101;
				18'b010101001110001100: oled_data = 16'b1101110011010101;
				18'b010101010000001100: oled_data = 16'b1101110011010101;
				18'b010101010010001100: oled_data = 16'b1101110011010101;
				18'b010101010100001100: oled_data = 16'b1101110011010101;
				18'b010101010110001100: oled_data = 16'b1101110010110101;
				18'b010101011000001100: oled_data = 16'b1101010001110100;
				18'b010101011010001100: oled_data = 16'b1101110011010110;
				18'b010101011100001100: oled_data = 16'b1101110011010101;
				18'b010101011110001100: oled_data = 16'b1101110011010101;
				18'b010101100000001100: oled_data = 16'b1101110011110110;
				18'b010101100010001100: oled_data = 16'b1101110011010101;
				18'b010101100100001100: oled_data = 16'b1101110011010101;
				18'b010101100110001100: oled_data = 16'b1101110011010110;
				18'b010101101000001100: oled_data = 16'b1110010011010110;
				18'b010101101010001100: oled_data = 16'b1101110011010101;
				18'b010101101100001100: oled_data = 16'b1101010010010101;
				18'b010101101110001100: oled_data = 16'b1101110011010101;
				18'b010101110000001100: oled_data = 16'b1101110011010101;
				18'b010101110010001100: oled_data = 16'b1101110011010101;
				18'b010101110100001100: oled_data = 16'b1101010010010101;
				18'b010101110110001100: oled_data = 16'b1101110011010101;
				18'b010101111000001100: oled_data = 16'b1101110011010101;
				18'b010101111010001100: oled_data = 16'b1101110011010110;
				18'b010101111100001100: oled_data = 16'b1101010010010101;
				18'b010101111110001100: oled_data = 16'b1101010010010100;
				18'b010110000000001100: oled_data = 16'b1101110011010101;
				18'b010110000010001100: oled_data = 16'b1101110011010101;
				18'b010110000100001100: oled_data = 16'b1101110010110101;
				18'b010110000110001100: oled_data = 16'b1101110101010111;
				18'b010110001000001100: oled_data = 16'b1111111100011101;
				18'b010110001010001100: oled_data = 16'b0111001101001101;
				18'b010110001100001100: oled_data = 16'b0001100100000100;
				18'b010110001110001100: oled_data = 16'b0010000101000101;
				18'b010110010000001100: oled_data = 16'b0010000101100110;
				18'b010110010010001100: oled_data = 16'b0010100101100110;
				18'b010110010100001100: oled_data = 16'b0010100110000111;
				18'b010110010110001100: oled_data = 16'b0010100110000111;
				18'b010110011000001100: oled_data = 16'b0010100110100111;
				18'b010110011010001100: oled_data = 16'b0110101010101010;
				18'b010110011100001100: oled_data = 16'b1011110001010001;
				18'b010110011110001100: oled_data = 16'b1110010011010100;
				18'b010110100000001100: oled_data = 16'b1101110000110001;
				18'b010110100010001100: oled_data = 16'b1100001100001100;
				18'b010110100100001100: oled_data = 16'b1010101001001001;
				18'b010110100110001100: oled_data = 16'b1010101000001000;
				18'b010100011000001101: oled_data = 16'b1001110001001100;
				18'b010100011010001101: oled_data = 16'b1000110010110000;
				18'b010100011100001101: oled_data = 16'b1000110100010010;
				18'b010100011110001101: oled_data = 16'b1010010111110111;
				18'b010100100000001101: oled_data = 16'b1011011000011000;
				18'b010100100010001101: oled_data = 16'b1100010100010110;
				18'b010100100100001101: oled_data = 16'b1101110011010110;
				18'b010100100110001101: oled_data = 16'b1110010011010110;
				18'b010100101000001101: oled_data = 16'b1101110011010101;
				18'b010100101010001101: oled_data = 16'b1101110011010101;
				18'b010100101100001101: oled_data = 16'b1101110011010101;
				18'b010100101110001101: oled_data = 16'b1101110011010101;
				18'b010100110000001101: oled_data = 16'b1101110011010110;
				18'b010100110010001101: oled_data = 16'b1101010010010101;
				18'b010100110100001101: oled_data = 16'b1101110010110101;
				18'b010100110110001101: oled_data = 16'b1101110011010110;
				18'b010100111000001101: oled_data = 16'b1101110011010101;
				18'b010100111010001101: oled_data = 16'b1110010011110110;
				18'b010100111100001101: oled_data = 16'b1110010011110110;
				18'b010100111110001101: oled_data = 16'b1101110011010101;
				18'b010101000000001101: oled_data = 16'b1101110011010101;
				18'b010101000010001101: oled_data = 16'b1101110011010101;
				18'b010101000100001101: oled_data = 16'b1101110011010101;
				18'b010101000110001101: oled_data = 16'b1101110011010101;
				18'b010101001000001101: oled_data = 16'b1101110011010101;
				18'b010101001010001101: oled_data = 16'b1101110011010101;
				18'b010101001100001101: oled_data = 16'b1101110011010101;
				18'b010101001110001101: oled_data = 16'b1101110011010101;
				18'b010101010000001101: oled_data = 16'b1101110011010101;
				18'b010101010010001101: oled_data = 16'b1101110011010101;
				18'b010101010100001101: oled_data = 16'b1101110011010101;
				18'b010101010110001101: oled_data = 16'b1101110010110101;
				18'b010101011000001101: oled_data = 16'b1101010010010101;
				18'b010101011010001101: oled_data = 16'b1101110011010110;
				18'b010101011100001101: oled_data = 16'b1101110011010101;
				18'b010101011110001101: oled_data = 16'b1101110011110110;
				18'b010101100000001101: oled_data = 16'b1110010101111000;
				18'b010101100010001101: oled_data = 16'b1101110011010101;
				18'b010101100100001101: oled_data = 16'b1101110011010101;
				18'b010101100110001101: oled_data = 16'b1101110011010101;
				18'b010101101000001101: oled_data = 16'b1101110011010101;
				18'b010101101010001101: oled_data = 16'b1101110011010101;
				18'b010101101100001101: oled_data = 16'b1101010010010100;
				18'b010101101110001101: oled_data = 16'b1101110011010101;
				18'b010101110000001101: oled_data = 16'b1101110011010101;
				18'b010101110010001101: oled_data = 16'b1101110011010110;
				18'b010101110100001101: oled_data = 16'b1101110010010101;
				18'b010101110110001101: oled_data = 16'b1101110011010101;
				18'b010101111000001101: oled_data = 16'b1101110011010101;
				18'b010101111010001101: oled_data = 16'b1101110011010101;
				18'b010101111100001101: oled_data = 16'b1101110010110101;
				18'b010101111110001101: oled_data = 16'b1101010010010100;
				18'b010110000000001101: oled_data = 16'b1101110011010101;
				18'b010110000010001101: oled_data = 16'b1101110011010101;
				18'b010110000100001101: oled_data = 16'b1101110010110101;
				18'b010110000110001101: oled_data = 16'b1101010011010101;
				18'b010110001000001101: oled_data = 16'b1111011011111100;
				18'b010110001010001101: oled_data = 16'b1010010011110100;
				18'b010110001100001101: oled_data = 16'b0001100100000100;
				18'b010110001110001101: oled_data = 16'b0010000101000101;
				18'b010110010000001101: oled_data = 16'b0010000101000110;
				18'b010110010010001101: oled_data = 16'b0010000101100110;
				18'b010110010100001101: oled_data = 16'b0010000101000110;
				18'b010110010110001101: oled_data = 16'b0100001000001000;
				18'b010110011000001101: oled_data = 16'b1010101111110000;
				18'b010110011010001101: oled_data = 16'b1110010100010100;
				18'b010110011100001101: oled_data = 16'b1110010010010010;
				18'b010110011110001101: oled_data = 16'b1100001100101101;
				18'b010110100000001101: oled_data = 16'b1011001001001001;
				18'b010110100010001101: oled_data = 16'b1011001000101000;
				18'b010110100100001101: oled_data = 16'b1010101000101000;
				18'b010110100110001101: oled_data = 16'b1010101000001000;
				18'b010100011000001110: oled_data = 16'b1001010011110001;
				18'b010100011010001110: oled_data = 16'b1000011000111001;
				18'b010100011100001110: oled_data = 16'b1010011100011100;
				18'b010100011110001110: oled_data = 16'b1010011011011011;
				18'b010100100000001110: oled_data = 16'b1001011010011010;
				18'b010100100010001110: oled_data = 16'b0111111000111001;
				18'b010100100100001110: oled_data = 16'b1000110110111000;
				18'b010100100110001110: oled_data = 16'b1011110100010110;
				18'b010100101000001110: oled_data = 16'b1110010010110110;
				18'b010100101010001110: oled_data = 16'b1101110011010110;
				18'b010100101100001110: oled_data = 16'b1101110011010101;
				18'b010100101110001110: oled_data = 16'b1101110011010101;
				18'b010100110000001110: oled_data = 16'b1101110010110101;
				18'b010100110010001110: oled_data = 16'b1101010001110100;
				18'b010100110100001110: oled_data = 16'b1101110011010110;
				18'b010100110110001110: oled_data = 16'b1101110011010101;
				18'b010100111000001110: oled_data = 16'b1101110011010110;
				18'b010100111010001110: oled_data = 16'b1110110100110111;
				18'b010100111100001110: oled_data = 16'b1110010011110110;
				18'b010100111110001110: oled_data = 16'b1101110011010101;
				18'b010101000000001110: oled_data = 16'b1101110011010101;
				18'b010101000010001110: oled_data = 16'b1101110011010101;
				18'b010101000100001110: oled_data = 16'b1101110011010101;
				18'b010101000110001110: oled_data = 16'b1101110010110101;
				18'b010101001000001110: oled_data = 16'b1101010010010100;
				18'b010101001010001110: oled_data = 16'b1101110011010101;
				18'b010101001100001110: oled_data = 16'b1101110011010101;
				18'b010101001110001110: oled_data = 16'b1101110011010101;
				18'b010101010000001110: oled_data = 16'b1101110011010101;
				18'b010101010010001110: oled_data = 16'b1101110011010101;
				18'b010101010100001110: oled_data = 16'b1101110011010101;
				18'b010101010110001110: oled_data = 16'b1101110010110101;
				18'b010101011000001110: oled_data = 16'b1101110010110101;
				18'b010101011010001110: oled_data = 16'b1101110011010110;
				18'b010101011100001110: oled_data = 16'b1101110011010101;
				18'b010101011110001110: oled_data = 16'b1110010011110110;
				18'b010101100000001110: oled_data = 16'b1110110110011000;
				18'b010101100010001110: oled_data = 16'b1101110011010101;
				18'b010101100100001110: oled_data = 16'b1101110011010101;
				18'b010101100110001110: oled_data = 16'b1101110011010101;
				18'b010101101000001110: oled_data = 16'b1101110011010101;
				18'b010101101010001110: oled_data = 16'b1101110011010110;
				18'b010101101100001110: oled_data = 16'b1101010001110100;
				18'b010101101110001110: oled_data = 16'b1101110011010101;
				18'b010101110000001110: oled_data = 16'b1101110011010101;
				18'b010101110010001110: oled_data = 16'b1101110011010110;
				18'b010101110100001110: oled_data = 16'b1101010010010101;
				18'b010101110110001110: oled_data = 16'b1101110010110101;
				18'b010101111000001110: oled_data = 16'b1101110011010110;
				18'b010101111010001110: oled_data = 16'b1101110011010110;
				18'b010101111100001110: oled_data = 16'b1101110011010101;
				18'b010101111110001110: oled_data = 16'b1101010001110100;
				18'b010110000000001110: oled_data = 16'b1101110011010101;
				18'b010110000010001110: oled_data = 16'b1101110011010101;
				18'b010110000100001110: oled_data = 16'b1101110010010101;
				18'b010110000110001110: oled_data = 16'b1101010010010100;
				18'b010110001000001110: oled_data = 16'b1110111001011010;
				18'b010110001010001110: oled_data = 16'b1100110111111000;
				18'b010110001100001110: oled_data = 16'b0010100101000101;
				18'b010110001110001110: oled_data = 16'b0010000100100101;
				18'b010110010000001110: oled_data = 16'b0010000100100101;
				18'b010110010010001110: oled_data = 16'b0010000100100101;
				18'b010110010100001110: oled_data = 16'b0110001010001010;
				18'b010110010110001110: oled_data = 16'b1101010010010010;
				18'b010110011000001110: oled_data = 16'b1110110011110100;
				18'b010110011010001110: oled_data = 16'b1101001111001111;
				18'b010110011100001110: oled_data = 16'b1011001010001010;
				18'b010110011110001110: oled_data = 16'b1011001000001000;
				18'b010110100000001110: oled_data = 16'b1011001000101001;
				18'b010110100010001110: oled_data = 16'b1011001000101000;
				18'b010110100100001110: oled_data = 16'b1010101000101000;
				18'b010110100110001110: oled_data = 16'b1010101000001000;
				18'b010100011000001111: oled_data = 16'b0111110110010110;
				18'b010100011010001111: oled_data = 16'b1000111010011011;
				18'b010100011100001111: oled_data = 16'b1011111100111100;
				18'b010100011110001111: oled_data = 16'b1011111100111101;
				18'b010100100000001111: oled_data = 16'b1011011100011100;
				18'b010100100010001111: oled_data = 16'b0111110111111001;
				18'b010100100100001111: oled_data = 16'b0111010111111010;
				18'b010100100110001111: oled_data = 16'b0111111000111010;
				18'b010100101000001111: oled_data = 16'b1011110100010111;
				18'b010100101010001111: oled_data = 16'b1110010011010101;
				18'b010100101100001111: oled_data = 16'b1101110011010101;
				18'b010100101110001111: oled_data = 16'b1101110011010101;
				18'b010100110000001111: oled_data = 16'b1101010001110100;
				18'b010100110010001111: oled_data = 16'b1101110010110101;
				18'b010100110100001111: oled_data = 16'b1101110011010101;
				18'b010100110110001111: oled_data = 16'b1101110011010101;
				18'b010100111000001111: oled_data = 16'b1110010011110110;
				18'b010100111010001111: oled_data = 16'b1110010011110110;
				18'b010100111100001111: oled_data = 16'b1101110011010101;
				18'b010100111110001111: oled_data = 16'b1101110011010101;
				18'b010101000000001111: oled_data = 16'b1101110011010101;
				18'b010101000010001111: oled_data = 16'b1101110011010101;
				18'b010101000100001111: oled_data = 16'b1101110011010101;
				18'b010101000110001111: oled_data = 16'b1101010010010100;
				18'b010101001000001111: oled_data = 16'b1101110010110101;
				18'b010101001010001111: oled_data = 16'b1101110011010101;
				18'b010101001100001111: oled_data = 16'b1101110011010101;
				18'b010101001110001111: oled_data = 16'b1101110010110101;
				18'b010101010000001111: oled_data = 16'b1101110010110101;
				18'b010101010010001111: oled_data = 16'b1101110011010101;
				18'b010101010100001111: oled_data = 16'b1101110011010110;
				18'b010101010110001111: oled_data = 16'b1101010010010100;
				18'b010101011000001111: oled_data = 16'b1101110010110101;
				18'b010101011010001111: oled_data = 16'b1101110011010101;
				18'b010101011100001111: oled_data = 16'b1101110011010101;
				18'b010101011110001111: oled_data = 16'b1110010100010110;
				18'b010101100000001111: oled_data = 16'b1110010110011000;
				18'b010101100010001111: oled_data = 16'b1101110011010101;
				18'b010101100100001111: oled_data = 16'b1101110011010101;
				18'b010101100110001111: oled_data = 16'b1101110011010101;
				18'b010101101000001111: oled_data = 16'b1101110011010101;
				18'b010101101010001111: oled_data = 16'b1101110011010110;
				18'b010101101100001111: oled_data = 16'b1101010001110100;
				18'b010101101110001111: oled_data = 16'b1101110010110101;
				18'b010101110000001111: oled_data = 16'b1101110011010101;
				18'b010101110010001111: oled_data = 16'b1101110011010110;
				18'b010101110100001111: oled_data = 16'b1101010010010100;
				18'b010101110110001111: oled_data = 16'b1101010010010101;
				18'b010101111000001111: oled_data = 16'b1101110011010110;
				18'b010101111010001111: oled_data = 16'b1101110011010110;
				18'b010101111100001111: oled_data = 16'b1101110011010101;
				18'b010101111110001111: oled_data = 16'b1101010001110100;
				18'b010110000000001111: oled_data = 16'b1101110011010101;
				18'b010110000010001111: oled_data = 16'b1101110011010101;
				18'b010110000100001111: oled_data = 16'b1101010001110100;
				18'b010110000110001111: oled_data = 16'b1101010001110100;
				18'b010110001000001111: oled_data = 16'b1110010110011000;
				18'b010110001010001111: oled_data = 16'b1110011010011010;
				18'b010110001100001111: oled_data = 16'b0100000110100111;
				18'b010110001110001111: oled_data = 16'b0010000100000101;
				18'b010110010000001111: oled_data = 16'b0010000100100101;
				18'b010110010010001111: oled_data = 16'b0111101100001100;
				18'b010110010100001111: oled_data = 16'b1110010100010100;
				18'b010110010110001111: oled_data = 16'b1110010010110010;
				18'b010110011000001111: oled_data = 16'b1100001100001100;
				18'b010110011010001111: oled_data = 16'b1011001000101001;
				18'b010110011100001111: oled_data = 16'b1011001000101001;
				18'b010110011110001111: oled_data = 16'b1011001000101001;
				18'b010110100000001111: oled_data = 16'b1011001000101001;
				18'b010110100010001111: oled_data = 16'b1011001000101000;
				18'b010110100100001111: oled_data = 16'b1010101000101000;
				18'b010110100110001111: oled_data = 16'b1010101000001000;
				18'b010100011000010000: oled_data = 16'b0110111000111001;
				18'b010100011010010000: oled_data = 16'b1000111010011011;
				18'b010100011100010000: oled_data = 16'b1011011100111100;
				18'b010100011110010000: oled_data = 16'b1001111001111010;
				18'b010100100000010000: oled_data = 16'b0111010101010111;
				18'b010100100010010000: oled_data = 16'b0100110001110101;
				18'b010100100100010000: oled_data = 16'b0101010010110110;
				18'b010100100110010000: oled_data = 16'b0110110111111010;
				18'b010100101000010000: oled_data = 16'b1001110101110111;
				18'b010100101010010000: oled_data = 16'b1110010010110101;
				18'b010100101100010000: oled_data = 16'b1101110011010101;
				18'b010100101110010000: oled_data = 16'b1101110010110101;
				18'b010100110000010000: oled_data = 16'b1101110010010101;
				18'b010100110010010000: oled_data = 16'b1101110011010110;
				18'b010100110100010000: oled_data = 16'b1101110011010101;
				18'b010100110110010000: oled_data = 16'b1101110011010101;
				18'b010100111000010000: oled_data = 16'b1101110011010110;
				18'b010100111010010000: oled_data = 16'b1101110011010110;
				18'b010100111100010000: oled_data = 16'b1101110011010101;
				18'b010100111110010000: oled_data = 16'b1101110011010101;
				18'b010101000000010000: oled_data = 16'b1101110011010101;
				18'b010101000010010000: oled_data = 16'b1101110011010101;
				18'b010101000100010000: oled_data = 16'b1101110010110101;
				18'b010101000110010000: oled_data = 16'b1101010010010101;
				18'b010101001000010000: oled_data = 16'b1101110011010110;
				18'b010101001010010000: oled_data = 16'b1101110011010101;
				18'b010101001100010000: oled_data = 16'b1101110011010110;
				18'b010101001110010000: oled_data = 16'b1101010010010100;
				18'b010101010000010000: oled_data = 16'b1101110010110101;
				18'b010101010010010000: oled_data = 16'b1101110011010101;
				18'b010101010100010000: oled_data = 16'b1101110011010110;
				18'b010101010110010000: oled_data = 16'b1101010010010100;
				18'b010101011000010000: oled_data = 16'b1101110010110101;
				18'b010101011010010000: oled_data = 16'b1101110011010101;
				18'b010101011100010000: oled_data = 16'b1101110011010101;
				18'b010101011110010000: oled_data = 16'b1110010011110110;
				18'b010101100000010000: oled_data = 16'b1110010100010110;
				18'b010101100010010000: oled_data = 16'b1101110011010101;
				18'b010101100100010000: oled_data = 16'b1101110011010101;
				18'b010101100110010000: oled_data = 16'b1101110011010101;
				18'b010101101000010000: oled_data = 16'b1101110011010101;
				18'b010101101010010000: oled_data = 16'b1101110011010110;
				18'b010101101100010000: oled_data = 16'b1101010010010100;
				18'b010101101110010000: oled_data = 16'b1101110010110101;
				18'b010101110000010000: oled_data = 16'b1101110011010101;
				18'b010101110010010000: oled_data = 16'b1101110011010110;
				18'b010101110100010000: oled_data = 16'b1101010010010100;
				18'b010101110110010000: oled_data = 16'b1101010001110100;
				18'b010101111000010000: oled_data = 16'b1101110011010110;
				18'b010101111010010000: oled_data = 16'b1101110011010110;
				18'b010101111100010000: oled_data = 16'b1101110011010101;
				18'b010101111110010000: oled_data = 16'b1101010010010100;
				18'b010110000000010000: oled_data = 16'b1101110011010110;
				18'b010110000010010000: oled_data = 16'b1101110011010110;
				18'b010110000100010000: oled_data = 16'b1101110010110101;
				18'b010110000110010000: oled_data = 16'b1101010001110100;
				18'b010110001000010000: oled_data = 16'b1101010100010110;
				18'b010110001010010000: oled_data = 16'b1111011011011011;
				18'b010110001100010000: oled_data = 16'b0100101000001000;
				18'b010110001110010000: oled_data = 16'b0010000100000100;
				18'b010110010000010000: oled_data = 16'b1000101100101101;
				18'b010110010010010000: oled_data = 16'b1110110100110101;
				18'b010110010100010000: oled_data = 16'b1101110001010001;
				18'b010110010110010000: oled_data = 16'b1011101010101010;
				18'b010110011000010000: oled_data = 16'b1011001000101001;
				18'b010110011010010000: oled_data = 16'b1011001000101001;
				18'b010110011100010000: oled_data = 16'b1011001001001001;
				18'b010110011110010000: oled_data = 16'b1011001000101001;
				18'b010110100000010000: oled_data = 16'b1011001000101001;
				18'b010110100010010000: oled_data = 16'b1011001000101000;
				18'b010110100100010000: oled_data = 16'b1010101000101000;
				18'b010110100110010000: oled_data = 16'b1010101000001000;
				18'b010100011000010001: oled_data = 16'b0111011000111010;
				18'b010100011010010001: oled_data = 16'b1000011000111001;
				18'b010100011100010001: oled_data = 16'b1001111001111010;
				18'b010100011110010001: oled_data = 16'b0100110001010100;
				18'b010100100000010001: oled_data = 16'b0100010001010101;
				18'b010100100010010001: oled_data = 16'b0100110001110110;
				18'b010100100100010001: oled_data = 16'b0100010001010110;
				18'b010100100110010001: oled_data = 16'b0110010101111001;
				18'b010100101000010001: oled_data = 16'b1001110101111000;
				18'b010100101010010001: oled_data = 16'b1110010010110110;
				18'b010100101100010001: oled_data = 16'b1101110011010101;
				18'b010100101110010001: oled_data = 16'b1101010010010100;
				18'b010100110000010001: oled_data = 16'b1101110011010110;
				18'b010100110010010001: oled_data = 16'b1101110011010101;
				18'b010100110100010001: oled_data = 16'b1101110011010101;
				18'b010100110110010001: oled_data = 16'b1101110011010101;
				18'b010100111000010001: oled_data = 16'b1101110011010101;
				18'b010100111010010001: oled_data = 16'b1101110011010101;
				18'b010100111100010001: oled_data = 16'b1101110011010101;
				18'b010100111110010001: oled_data = 16'b1101110011010101;
				18'b010101000000010001: oled_data = 16'b1101110011010101;
				18'b010101000010010001: oled_data = 16'b1101110011010110;
				18'b010101000100010001: oled_data = 16'b1101010001110100;
				18'b010101000110010001: oled_data = 16'b1101110010110101;
				18'b010101001000010001: oled_data = 16'b1101110011010101;
				18'b010101001010010001: oled_data = 16'b1101110011010101;
				18'b010101001100010001: oled_data = 16'b1101110011010110;
				18'b010101001110010001: oled_data = 16'b1101010001110100;
				18'b010101010000010001: oled_data = 16'b1101110010110101;
				18'b010101010010010001: oled_data = 16'b1101110011010101;
				18'b010101010100010001: oled_data = 16'b1101110011010101;
				18'b010101010110010001: oled_data = 16'b1101010010010100;
				18'b010101011000010001: oled_data = 16'b1101110011010101;
				18'b010101011010010001: oled_data = 16'b1101110011010101;
				18'b010101011100010001: oled_data = 16'b1101110011010101;
				18'b010101011110010001: oled_data = 16'b1101110011010101;
				18'b010101100000010001: oled_data = 16'b1101110011010101;
				18'b010101100010010001: oled_data = 16'b1101110011010101;
				18'b010101100100010001: oled_data = 16'b1101110011010101;
				18'b010101100110010001: oled_data = 16'b1101110011010101;
				18'b010101101000010001: oled_data = 16'b1101110011010101;
				18'b010101101010010001: oled_data = 16'b1101110011010110;
				18'b010101101100010001: oled_data = 16'b1101010010010100;
				18'b010101101110010001: oled_data = 16'b1101110010110101;
				18'b010101110000010001: oled_data = 16'b1101110011010101;
				18'b010101110010010001: oled_data = 16'b1101110011010110;
				18'b010101110100010001: oled_data = 16'b1101010010010101;
				18'b010101110110010001: oled_data = 16'b1101010001110100;
				18'b010101111000010001: oled_data = 16'b1110010011010110;
				18'b010101111010010001: oled_data = 16'b1101110011010110;
				18'b010101111100010001: oled_data = 16'b1101110011010110;
				18'b010101111110010001: oled_data = 16'b1100110000110011;
				18'b010110000000010001: oled_data = 16'b1101110011010110;
				18'b010110000010010001: oled_data = 16'b1110010011010110;
				18'b010110000100010001: oled_data = 16'b1101110011010101;
				18'b010110000110010001: oled_data = 16'b1101010001110100;
				18'b010110001000010001: oled_data = 16'b1100110011010101;
				18'b010110001010010001: oled_data = 16'b1111011011011100;
				18'b010110001100010001: oled_data = 16'b0101101010001011;
				18'b010110001110010001: oled_data = 16'b1000101100101101;
				18'b010110010000010001: oled_data = 16'b1110110100010101;
				18'b010110010010010001: oled_data = 16'b1101010000010000;
				18'b010110010100010001: oled_data = 16'b1011001001101010;
				18'b010110010110010001: oled_data = 16'b1011001000101001;
				18'b010110011000010001: oled_data = 16'b1011001001001001;
				18'b010110011010010001: oled_data = 16'b1011001000101001;
				18'b010110011100010001: oled_data = 16'b1011001001001001;
				18'b010110011110010001: oled_data = 16'b1011001000101001;
				18'b010110100000010001: oled_data = 16'b1011001000101001;
				18'b010110100010010001: oled_data = 16'b1011001000101000;
				18'b010110100100010001: oled_data = 16'b1011001000001000;
				18'b010110100110010001: oled_data = 16'b1011001000001000;
				18'b010100011000010010: oled_data = 16'b0110111000011001;
				18'b010100011010010010: oled_data = 16'b0110110101111000;
				18'b010100011100010010: oled_data = 16'b0111010101011000;
				18'b010100011110010010: oled_data = 16'b0100010000110101;
				18'b010100100000010010: oled_data = 16'b0100010001110101;
				18'b010100100010010010: oled_data = 16'b0100110001110101;
				18'b010100100100010010: oled_data = 16'b0100110001010101;
				18'b010100100110010010: oled_data = 16'b0101110101011000;
				18'b010100101000010010: oled_data = 16'b1010010101010111;
				18'b010100101010010010: oled_data = 16'b1110010011010110;
				18'b010100101100010010: oled_data = 16'b1101110010110101;
				18'b010100101110010010: oled_data = 16'b1101110010110101;
				18'b010100110000010010: oled_data = 16'b1101110011010101;
				18'b010100110010010010: oled_data = 16'b1101110011010110;
				18'b010100110100010010: oled_data = 16'b1101010010010101;
				18'b010100110110010010: oled_data = 16'b1101010010010101;
				18'b010100111000010010: oled_data = 16'b1101110011010110;
				18'b010100111010010010: oled_data = 16'b1101110011010101;
				18'b010100111100010010: oled_data = 16'b1101110011010101;
				18'b010100111110010010: oled_data = 16'b1101110011010101;
				18'b010101000000010010: oled_data = 16'b1101110011010101;
				18'b010101000010010010: oled_data = 16'b1101110011010101;
				18'b010101000100010010: oled_data = 16'b1101010010010100;
				18'b010101000110010010: oled_data = 16'b1101110011010101;
				18'b010101001000010010: oled_data = 16'b1101110011010101;
				18'b010101001010010010: oled_data = 16'b1101110011010101;
				18'b010101001100010010: oled_data = 16'b1101110011010101;
				18'b010101001110010010: oled_data = 16'b1101010001110100;
				18'b010101010000010010: oled_data = 16'b1101110011010101;
				18'b010101010010010010: oled_data = 16'b1101110011010101;
				18'b010101010100010010: oled_data = 16'b1101110011010101;
				18'b010101010110010010: oled_data = 16'b1101110010010101;
				18'b010101011000010010: oled_data = 16'b1110010011110110;
				18'b010101011010010010: oled_data = 16'b1110010011010110;
				18'b010101011100010010: oled_data = 16'b1101110011010101;
				18'b010101011110010010: oled_data = 16'b1101110011010101;
				18'b010101100000010010: oled_data = 16'b1101110011010101;
				18'b010101100010010010: oled_data = 16'b1101110011010101;
				18'b010101100100010010: oled_data = 16'b1101110011010101;
				18'b010101100110010010: oled_data = 16'b1101110011010101;
				18'b010101101000010010: oled_data = 16'b1101110011010101;
				18'b010101101010010010: oled_data = 16'b1101110011010110;
				18'b010101101100010010: oled_data = 16'b1101010001110100;
				18'b010101101110010010: oled_data = 16'b1101110010110101;
				18'b010101110000010010: oled_data = 16'b1101110011010101;
				18'b010101110010010010: oled_data = 16'b1101110011010110;
				18'b010101110100010010: oled_data = 16'b1101110010110101;
				18'b010101110110010010: oled_data = 16'b1101010010010100;
				18'b010101111000010010: oled_data = 16'b1101110011010110;
				18'b010101111010010010: oled_data = 16'b1101110011010110;
				18'b010101111100010010: oled_data = 16'b1101110011010110;
				18'b010101111110010010: oled_data = 16'b1100001111110010;
				18'b010110000000010010: oled_data = 16'b1101110011010101;
				18'b010110000010010010: oled_data = 16'b1110010011010110;
				18'b010110000100010010: oled_data = 16'b1101110011010110;
				18'b010110000110010010: oled_data = 16'b1101010001110100;
				18'b010110001000010010: oled_data = 16'b1101010011010101;
				18'b010110001010010010: oled_data = 16'b1110111001011010;
				18'b010110001100010010: oled_data = 16'b1011010000110010;
				18'b010110001110010010: oled_data = 16'b1110010011110100;
				18'b010110010000010010: oled_data = 16'b1101110000110000;
				18'b010110010010010010: oled_data = 16'b1011001001101001;
				18'b010110010100010010: oled_data = 16'b1011001001001001;
				18'b010110010110010010: oled_data = 16'b1011001001001001;
				18'b010110011000010010: oled_data = 16'b1011001001001001;
				18'b010110011010010010: oled_data = 16'b1011001000101001;
				18'b010110011100010010: oled_data = 16'b1011001001001001;
				18'b010110011110010010: oled_data = 16'b1011001000101001;
				18'b010110100000010010: oled_data = 16'b1011001000101001;
				18'b010110100010010010: oled_data = 16'b1011001000101000;
				18'b010110100100010010: oled_data = 16'b1011001000101000;
				18'b010110100110010010: oled_data = 16'b1011001000001000;
				18'b010100011000010011: oled_data = 16'b0110110111111001;
				18'b010100011010010011: oled_data = 16'b0101010011010110;
				18'b010100011100010011: oled_data = 16'b0101010011010111;
				18'b010100011110010011: oled_data = 16'b0100110001010101;
				18'b010100100000010011: oled_data = 16'b0100010001110101;
				18'b010100100010010011: oled_data = 16'b0100010001110101;
				18'b010100100100010011: oled_data = 16'b0100010001010101;
				18'b010100100110010011: oled_data = 16'b0101110101010111;
				18'b010100101000010011: oled_data = 16'b1011010100110110;
				18'b010100101010010011: oled_data = 16'b1110010010110101;
				18'b010100101100010011: oled_data = 16'b1101010001110100;
				18'b010100101110010011: oled_data = 16'b1101110011010110;
				18'b010100110000010011: oled_data = 16'b1101110011010101;
				18'b010100110010010011: oled_data = 16'b1101110011010101;
				18'b010100110100010011: oled_data = 16'b1100010000010010;
				18'b010100110110010011: oled_data = 16'b1101110010110101;
				18'b010100111000010011: oled_data = 16'b1101110011010101;
				18'b010100111010010011: oled_data = 16'b1101110011010101;
				18'b010100111100010011: oled_data = 16'b1101110011010101;
				18'b010100111110010011: oled_data = 16'b1101110011010101;
				18'b010101000000010011: oled_data = 16'b1101110011010110;
				18'b010101000010010011: oled_data = 16'b1101010010010101;
				18'b010101000100010011: oled_data = 16'b1101010010010101;
				18'b010101000110010011: oled_data = 16'b1101110011010101;
				18'b010101001000010011: oled_data = 16'b1101110011010101;
				18'b010101001010010011: oled_data = 16'b1101110011010101;
				18'b010101001100010011: oled_data = 16'b1101110010110101;
				18'b010101001110010011: oled_data = 16'b1100110000110011;
				18'b010101010000010011: oled_data = 16'b1101110011010110;
				18'b010101010010010011: oled_data = 16'b1101110011010101;
				18'b010101010100010011: oled_data = 16'b1101110011010101;
				18'b010101010110010011: oled_data = 16'b1101010001110100;
				18'b010101011000010011: oled_data = 16'b1110010011010110;
				18'b010101011010010011: oled_data = 16'b1110010011110110;
				18'b010101011100010011: oled_data = 16'b1101110011010110;
				18'b010101011110010011: oled_data = 16'b1101110011010101;
				18'b010101100000010011: oled_data = 16'b1101110011010101;
				18'b010101100010010011: oled_data = 16'b1101110011010101;
				18'b010101100100010011: oled_data = 16'b1101110011010101;
				18'b010101100110010011: oled_data = 16'b1101110011010101;
				18'b010101101000010011: oled_data = 16'b1101110011010101;
				18'b010101101010010011: oled_data = 16'b1101110011010110;
				18'b010101101100010011: oled_data = 16'b1101010001110100;
				18'b010101101110010011: oled_data = 16'b1101110010110101;
				18'b010101110000010011: oled_data = 16'b1101110011010101;
				18'b010101110010010011: oled_data = 16'b1101110011010110;
				18'b010101110100010011: oled_data = 16'b1101010010010100;
				18'b010101110110010011: oled_data = 16'b1100010001110011;
				18'b010101111000010011: oled_data = 16'b1101110011010110;
				18'b010101111010010011: oled_data = 16'b1101110011010110;
				18'b010101111100010011: oled_data = 16'b1101110011010110;
				18'b010101111110010011: oled_data = 16'b1011101110110001;
				18'b010110000000010011: oled_data = 16'b1101110010110101;
				18'b010110000010010011: oled_data = 16'b1110010011110110;
				18'b010110000100010011: oled_data = 16'b1101110011010110;
				18'b010110000110010011: oled_data = 16'b1101010001110100;
				18'b010110001000010011: oled_data = 16'b1101110010110101;
				18'b010110001010010011: oled_data = 16'b1101110100010110;
				18'b010110001100010011: oled_data = 16'b1110010100010100;
				18'b010110001110010011: oled_data = 16'b1101110001010001;
				18'b010110010000010011: oled_data = 16'b1011001010001010;
				18'b010110010010010011: oled_data = 16'b1011001001001001;
				18'b010110010100010011: oled_data = 16'b1011001001001001;
				18'b010110010110010011: oled_data = 16'b1011001001001001;
				18'b010110011000010011: oled_data = 16'b1011001001001001;
				18'b010110011010010011: oled_data = 16'b1011001000101001;
				18'b010110011100010011: oled_data = 16'b1011001001001001;
				18'b010110011110010011: oled_data = 16'b1011001000101001;
				18'b010110100000010011: oled_data = 16'b1011001000101001;
				18'b010110100010010011: oled_data = 16'b1011001000101001;
				18'b010110100100010011: oled_data = 16'b1011001000101000;
				18'b010110100110010011: oled_data = 16'b1011001000001000;
				18'b010100011000010100: oled_data = 16'b0110110111111001;
				18'b010100011010010100: oled_data = 16'b0100010010010101;
				18'b010100011100010100: oled_data = 16'b0100110001110110;
				18'b010100011110010100: oled_data = 16'b0100110001010110;
				18'b010100100000010100: oled_data = 16'b0100010001010101;
				18'b010100100010010100: oled_data = 16'b0100010001110101;
				18'b010100100100010100: oled_data = 16'b0100010001110101;
				18'b010100100110010100: oled_data = 16'b0110110100110111;
				18'b010100101000010100: oled_data = 16'b1100110011010110;
				18'b010100101010010100: oled_data = 16'b1101110010010101;
				18'b010100101100010100: oled_data = 16'b1101010010010101;
				18'b010100101110010100: oled_data = 16'b1101110011010110;
				18'b010100110000010100: oled_data = 16'b1101110011010101;
				18'b010100110010010100: oled_data = 16'b1101010010010100;
				18'b010100110100010100: oled_data = 16'b1100110000110011;
				18'b010100110110010100: oled_data = 16'b1101110011010110;
				18'b010100111000010100: oled_data = 16'b1101110011010101;
				18'b010100111010010100: oled_data = 16'b1101110011010101;
				18'b010100111100010100: oled_data = 16'b1101110011010101;
				18'b010100111110010100: oled_data = 16'b1101110011010101;
				18'b010101000000010100: oled_data = 16'b1101110011010110;
				18'b010101000010010100: oled_data = 16'b1101010001110100;
				18'b010101000100010100: oled_data = 16'b1101110010110101;
				18'b010101000110010100: oled_data = 16'b1101110011010101;
				18'b010101001000010100: oled_data = 16'b1101110011010101;
				18'b010101001010010100: oled_data = 16'b1110010011010110;
				18'b010101001100010100: oled_data = 16'b1101010010010100;
				18'b010101001110010100: oled_data = 16'b1101010001110100;
				18'b010101010000010100: oled_data = 16'b1101110011010110;
				18'b010101010010010100: oled_data = 16'b1101110011010101;
				18'b010101010100010100: oled_data = 16'b1101110010110101;
				18'b010101010110010100: oled_data = 16'b1100110000110011;
				18'b010101011000010100: oled_data = 16'b1101110011010110;
				18'b010101011010010100: oled_data = 16'b1101110011010110;
				18'b010101011100010100: oled_data = 16'b1101110011010101;
				18'b010101011110010100: oled_data = 16'b1101110011010101;
				18'b010101100000010100: oled_data = 16'b1101110011010101;
				18'b010101100010010100: oled_data = 16'b1101110011010101;
				18'b010101100100010100: oled_data = 16'b1101110011010101;
				18'b010101100110010100: oled_data = 16'b1101110011010101;
				18'b010101101000010100: oled_data = 16'b1101110011010101;
				18'b010101101010010100: oled_data = 16'b1101110011010110;
				18'b010101101100010100: oled_data = 16'b1101010001110100;
				18'b010101101110010100: oled_data = 16'b1101110010110101;
				18'b010101110000010100: oled_data = 16'b1101110011010101;
				18'b010101110010010100: oled_data = 16'b1101110011010101;
				18'b010101110100010100: oled_data = 16'b1101010010110101;
				18'b010101110110010100: oled_data = 16'b1100110001110100;
				18'b010101111000010100: oled_data = 16'b1101110011010110;
				18'b010101111010010100: oled_data = 16'b1101110011010110;
				18'b010101111100010100: oled_data = 16'b1101110010110110;
				18'b010101111110010100: oled_data = 16'b1011101110010001;
				18'b010110000000010100: oled_data = 16'b1101110010010101;
				18'b010110000010010100: oled_data = 16'b1110010011110110;
				18'b010110000100010100: oled_data = 16'b1101110011010110;
				18'b010110000110010100: oled_data = 16'b1101110010010101;
				18'b010110001000010100: oled_data = 16'b1101010010010100;
				18'b010110001010010100: oled_data = 16'b1110010011010101;
				18'b010110001100010100: oled_data = 16'b1110010011010011;
				18'b010110001110010100: oled_data = 16'b1011101011001011;
				18'b010110010000010100: oled_data = 16'b1011001001001001;
				18'b010110010010010100: oled_data = 16'b1011101001001001;
				18'b010110010100010100: oled_data = 16'b1011001001001001;
				18'b010110010110010100: oled_data = 16'b1011001001001001;
				18'b010110011000010100: oled_data = 16'b1011001001001001;
				18'b010110011010010100: oled_data = 16'b1011001000101001;
				18'b010110011100010100: oled_data = 16'b1011001001001001;
				18'b010110011110010100: oled_data = 16'b1011001000101001;
				18'b010110100000010100: oled_data = 16'b1010101000001000;
				18'b010110100010010100: oled_data = 16'b1011001000101001;
				18'b010110100100010100: oled_data = 16'b1011001000101000;
				18'b010110100110010100: oled_data = 16'b1011001000001000;
				18'b010100011000010101: oled_data = 16'b0111010110111001;
				18'b010100011010010101: oled_data = 16'b0100110010010110;
				18'b010100011100010101: oled_data = 16'b0100110001010110;
				18'b010100011110010101: oled_data = 16'b0100110001010110;
				18'b010100100000010101: oled_data = 16'b0100110001010101;
				18'b010100100010010101: oled_data = 16'b0100010001010101;
				18'b010100100100010101: oled_data = 16'b0100110010010110;
				18'b010100100110010101: oled_data = 16'b1000110100010110;
				18'b010100101000010101: oled_data = 16'b1101010010110101;
				18'b010100101010010101: oled_data = 16'b1101010001110100;
				18'b010100101100010101: oled_data = 16'b1101110011010110;
				18'b010100101110010101: oled_data = 16'b1101110011010101;
				18'b010100110000010101: oled_data = 16'b1101110011010101;
				18'b010100110010010101: oled_data = 16'b1101010001110100;
				18'b010100110100010101: oled_data = 16'b1101010010010100;
				18'b010100110110010101: oled_data = 16'b1101110011010110;
				18'b010100111000010101: oled_data = 16'b1101110011010101;
				18'b010100111010010101: oled_data = 16'b1101110011010101;
				18'b010100111100010101: oled_data = 16'b1101110011010101;
				18'b010100111110010101: oled_data = 16'b1101110011010101;
				18'b010101000000010101: oled_data = 16'b1101110011010101;
				18'b010101000010010101: oled_data = 16'b1101010001110100;
				18'b010101000100010101: oled_data = 16'b1101110011010101;
				18'b010101000110010101: oled_data = 16'b1101110011010101;
				18'b010101001000010101: oled_data = 16'b1101110011010101;
				18'b010101001010010101: oled_data = 16'b1110010011010110;
				18'b010101001100010101: oled_data = 16'b1101010001110100;
				18'b010101001110010101: oled_data = 16'b1101010010010100;
				18'b010101010000010101: oled_data = 16'b1101110011010110;
				18'b010101010010010101: oled_data = 16'b1101110011010110;
				18'b010101010100010101: oled_data = 16'b1101110010010101;
				18'b010101010110010101: oled_data = 16'b1101010001110100;
				18'b010101011000010101: oled_data = 16'b1101110011010110;
				18'b010101011010010101: oled_data = 16'b1101110011010101;
				18'b010101011100010101: oled_data = 16'b1101110010110101;
				18'b010101011110010101: oled_data = 16'b1101110011010101;
				18'b010101100000010101: oled_data = 16'b1110010011010110;
				18'b010101100010010101: oled_data = 16'b1110010011010110;
				18'b010101100100010101: oled_data = 16'b1101110011010101;
				18'b010101100110010101: oled_data = 16'b1101110011010101;
				18'b010101101000010101: oled_data = 16'b1101110010110101;
				18'b010101101010010101: oled_data = 16'b1101110011010101;
				18'b010101101100010101: oled_data = 16'b1101010001110100;
				18'b010101101110010101: oled_data = 16'b1101110010110101;
				18'b010101110000010101: oled_data = 16'b1101110010110101;
				18'b010101110010010101: oled_data = 16'b1101010010110101;
				18'b010101110100010101: oled_data = 16'b1100110010110101;
				18'b010101110110010101: oled_data = 16'b1100110010010101;
				18'b010101111000010101: oled_data = 16'b1101110011010110;
				18'b010101111010010101: oled_data = 16'b1101110011010110;
				18'b010101111100010101: oled_data = 16'b1101110010110101;
				18'b010101111110010101: oled_data = 16'b1011001101110000;
				18'b010110000000010101: oled_data = 16'b1101010001110100;
				18'b010110000010010101: oled_data = 16'b1101110011010110;
				18'b010110000100010101: oled_data = 16'b1101110011010110;
				18'b010110000110010101: oled_data = 16'b1101010010010100;
				18'b010110001000010101: oled_data = 16'b1101110010110011;
				18'b010110001010010101: oled_data = 16'b1110110011110100;
				18'b010110001100010101: oled_data = 16'b1100001100101101;
				18'b010110001110010101: oled_data = 16'b1011001000101001;
				18'b010110010000010101: oled_data = 16'b1011101001001001;
				18'b010110010010010101: oled_data = 16'b1011101000101001;
				18'b010110010100010101: oled_data = 16'b1011001001001001;
				18'b010110010110010101: oled_data = 16'b1011001001001001;
				18'b010110011000010101: oled_data = 16'b1011001001001001;
				18'b010110011010010101: oled_data = 16'b1011001001001001;
				18'b010110011100010101: oled_data = 16'b1011001000101001;
				18'b010110011110010101: oled_data = 16'b1010001000001000;
				18'b010110100000010101: oled_data = 16'b1010101000001000;
				18'b010110100010010101: oled_data = 16'b1011001000101001;
				18'b010110100100010101: oled_data = 16'b1011001000101000;
				18'b010110100110010101: oled_data = 16'b1011001000001000;
				18'b010100011000010110: oled_data = 16'b1011010010110100;
				18'b010100011010010110: oled_data = 16'b0111110001110110;
				18'b010100011100010110: oled_data = 16'b0100110001110110;
				18'b010100011110010110: oled_data = 16'b0100110001110101;
				18'b010100100000010110: oled_data = 16'b0100110001010101;
				18'b010100100010010110: oled_data = 16'b0100110001110101;
				18'b010100100100010110: oled_data = 16'b0110010100111000;
				18'b010100100110010110: oled_data = 16'b1010010010110110;
				18'b010100101000010110: oled_data = 16'b1101110010110101;
				18'b010100101010010110: oled_data = 16'b1101110010010101;
				18'b010100101100010110: oled_data = 16'b1101110011010110;
				18'b010100101110010110: oled_data = 16'b1101110011010101;
				18'b010100110000010110: oled_data = 16'b1101110010110101;
				18'b010100110010010110: oled_data = 16'b1101010001110100;
				18'b010100110100010110: oled_data = 16'b1101110010110101;
				18'b010100110110010110: oled_data = 16'b1101110011010101;
				18'b010100111000010110: oled_data = 16'b1101110011010101;
				18'b010100111010010110: oled_data = 16'b1101110011010101;
				18'b010100111100010110: oled_data = 16'b1101110011010101;
				18'b010100111110010110: oled_data = 16'b1101110011010101;
				18'b010101000000010110: oled_data = 16'b1101110011010101;
				18'b010101000010010110: oled_data = 16'b1101110010010101;
				18'b010101000100010110: oled_data = 16'b1110010011010101;
				18'b010101000110010110: oled_data = 16'b1110010011010101;
				18'b010101001000010110: oled_data = 16'b1110010011010101;
				18'b010101001010010110: oled_data = 16'b1101110011010101;
				18'b010101001100010110: oled_data = 16'b1101010010010100;
				18'b010101001110010110: oled_data = 16'b1101110010110101;
				18'b010101010000010110: oled_data = 16'b1101110011010101;
				18'b010101010010010110: oled_data = 16'b1101110011010110;
				18'b010101010100010110: oled_data = 16'b1101010010010100;
				18'b010101010110010110: oled_data = 16'b1101010010010100;
				18'b010101011000010110: oled_data = 16'b1101110011010110;
				18'b010101011010010110: oled_data = 16'b1101110011010101;
				18'b010101011100010110: oled_data = 16'b1101110010110101;
				18'b010101011110010110: oled_data = 16'b1110010011010101;
				18'b010101100000010110: oled_data = 16'b1110010011010110;
				18'b010101100010010110: oled_data = 16'b1110010011010110;
				18'b010101100100010110: oled_data = 16'b1110010011010110;
				18'b010101100110010110: oled_data = 16'b1110010011010110;
				18'b010101101000010110: oled_data = 16'b1101010010010100;
				18'b010101101010010110: oled_data = 16'b1101110011010101;
				18'b010101101100010110: oled_data = 16'b1101010001110100;
				18'b010101101110010110: oled_data = 16'b1101010001110100;
				18'b010101110000010110: oled_data = 16'b1101110011010101;
				18'b010101110010010110: oled_data = 16'b1011110000010010;
				18'b010101110100010110: oled_data = 16'b1000001010001011;
				18'b010101110110010110: oled_data = 16'b1100110010010100;
				18'b010101111000010110: oled_data = 16'b1110010011010110;
				18'b010101111010010110: oled_data = 16'b1101110011010110;
				18'b010101111100010110: oled_data = 16'b1101010001110100;
				18'b010101111110010110: oled_data = 16'b1011001101110000;
				18'b010110000000010110: oled_data = 16'b1101010001010100;
				18'b010110000010010110: oled_data = 16'b1110010011010110;
				18'b010110000100010110: oled_data = 16'b1101110011010101;
				18'b010110000110010110: oled_data = 16'b1101010010010100;
				18'b010110001000010110: oled_data = 16'b1110110100010100;
				18'b010110001010010110: oled_data = 16'b1101010000010000;
				18'b010110001100010110: oled_data = 16'b1011001001001001;
				18'b010110001110010110: oled_data = 16'b1011101001001001;
				18'b010110010000010110: oled_data = 16'b1011101001001001;
				18'b010110010010010110: oled_data = 16'b1011101001001001;
				18'b010110010100010110: oled_data = 16'b1011001001001001;
				18'b010110010110010110: oled_data = 16'b1011001001001001;
				18'b010110011000010110: oled_data = 16'b1011001001001001;
				18'b010110011010010110: oled_data = 16'b1010101000101000;
				18'b010110011100010110: oled_data = 16'b1010001000001000;
				18'b010110011110010110: oled_data = 16'b1011001000101001;
				18'b010110100000010110: oled_data = 16'b1011001000101001;
				18'b010110100010010110: oled_data = 16'b1011001000101001;
				18'b010110100100010110: oled_data = 16'b1011001000101000;
				18'b010110100110010110: oled_data = 16'b1011001000001000;
				18'b010100011000010111: oled_data = 16'b1101011001010000;
				18'b010100011010010111: oled_data = 16'b1011010111010000;
				18'b010100011100010111: oled_data = 16'b1001010110110101;
				18'b010100011110010111: oled_data = 16'b0111010110010111;
				18'b010100100000010111: oled_data = 16'b0110110101111001;
				18'b010100100010010111: oled_data = 16'b0110110110111010;
				18'b010100100100010111: oled_data = 16'b0111110101011000;
				18'b010100100110010111: oled_data = 16'b1100110001010101;
				18'b010100101000010111: oled_data = 16'b1101010010010101;
				18'b010100101010010111: oled_data = 16'b1101110010110101;
				18'b010100101100010111: oled_data = 16'b1101110011010101;
				18'b010100101110010111: oled_data = 16'b1101110011010101;
				18'b010100110000010111: oled_data = 16'b1101010010010100;
				18'b010100110010010111: oled_data = 16'b1101010010010100;
				18'b010100110100010111: oled_data = 16'b1101110010110101;
				18'b010100110110010111: oled_data = 16'b1101110011010101;
				18'b010100111000010111: oled_data = 16'b1101110011010101;
				18'b010100111010010111: oled_data = 16'b1101110011010101;
				18'b010100111100010111: oled_data = 16'b1101110011010101;
				18'b010100111110010111: oled_data = 16'b1101110011010110;
				18'b010101000000010111: oled_data = 16'b1101010010010101;
				18'b010101000010010111: oled_data = 16'b1101110010110101;
				18'b010101000100010111: oled_data = 16'b1101110011010110;
				18'b010101000110010111: oled_data = 16'b1101110011010101;
				18'b010101001000010111: oled_data = 16'b1101110011010110;
				18'b010101001010010111: oled_data = 16'b1101010011010101;
				18'b010101001100010111: oled_data = 16'b1100010011010100;
				18'b010101001110010111: oled_data = 16'b1101110010110101;
				18'b010101010000010111: oled_data = 16'b1101110011010101;
				18'b010101010010010111: oled_data = 16'b1101110011010101;
				18'b010101010100010111: oled_data = 16'b1101010010110100;
				18'b010101010110010111: oled_data = 16'b1101010011010101;
				18'b010101011000010111: oled_data = 16'b1110010011010110;
				18'b010101011010010111: oled_data = 16'b1101110011010101;
				18'b010101011100010111: oled_data = 16'b1110010011010101;
				18'b010101011110010111: oled_data = 16'b1101110011010110;
				18'b010101100000010111: oled_data = 16'b1110010011010110;
				18'b010101100010010111: oled_data = 16'b1101110011010110;
				18'b010101100100010111: oled_data = 16'b1101110011010101;
				18'b010101100110010111: oled_data = 16'b1101110011010110;
				18'b010101101000010111: oled_data = 16'b1101010010010100;
				18'b010101101010010111: oled_data = 16'b1101110011110101;
				18'b010101101100010111: oled_data = 16'b1100010000110011;
				18'b010101101110010111: oled_data = 16'b1101010001110100;
				18'b010101110000010111: oled_data = 16'b1110010100010110;
				18'b010101110010010111: oled_data = 16'b1000001011001100;
				18'b010101110100010111: oled_data = 16'b0111001011101100;
				18'b010101110110010111: oled_data = 16'b1101010100010110;
				18'b010101111000010111: oled_data = 16'b1101110011010110;
				18'b010101111010010111: oled_data = 16'b1110010011010110;
				18'b010101111100010111: oled_data = 16'b1100001111110010;
				18'b010101111110010111: oled_data = 16'b1011001101110000;
				18'b010110000000010111: oled_data = 16'b1100110001010100;
				18'b010110000010010111: oled_data = 16'b1101110011110110;
				18'b010110000100010111: oled_data = 16'b1101010001110011;
				18'b010110000110010111: oled_data = 16'b1110010011110100;
				18'b010110001000010111: oled_data = 16'b1110010010110010;
				18'b010110001010010111: oled_data = 16'b1011101010101010;
				18'b010110001100010111: oled_data = 16'b1011001001001001;
				18'b010110001110010111: oled_data = 16'b1011001001001001;
				18'b010110010000010111: oled_data = 16'b1011001001001001;
				18'b010110010010010111: oled_data = 16'b1011001001001001;
				18'b010110010100010111: oled_data = 16'b1011001001001001;
				18'b010110010110010111: oled_data = 16'b1011001001001001;
				18'b010110011000010111: oled_data = 16'b1011001000101001;
				18'b010110011010010111: oled_data = 16'b1010001000001000;
				18'b010110011100010111: oled_data = 16'b1011001001001001;
				18'b010110011110010111: oled_data = 16'b1011001000101001;
				18'b010110100000010111: oled_data = 16'b1011001000101001;
				18'b010110100010010111: oled_data = 16'b1011001000101001;
				18'b010110100100010111: oled_data = 16'b1011001000101000;
				18'b010110100110010111: oled_data = 16'b1011001000001000;
				18'b010100011000011000: oled_data = 16'b1110111100010101;
				18'b010100011010011000: oled_data = 16'b1101111001110001;
				18'b010100011100011000: oled_data = 16'b1011110101101011;
				18'b010100011110011000: oled_data = 16'b1011010101101101;
				18'b010100100000011000: oled_data = 16'b1011010111010001;
				18'b010100100010011000: oled_data = 16'b1010110111110011;
				18'b010100100100011000: oled_data = 16'b1010010001010010;
				18'b010100100110011000: oled_data = 16'b1101010001110101;
				18'b010100101000011000: oled_data = 16'b1101010010010101;
				18'b010100101010011000: oled_data = 16'b1101110011010110;
				18'b010100101100011000: oled_data = 16'b1101110011010101;
				18'b010100101110011000: oled_data = 16'b1101010010010101;
				18'b010100110000011000: oled_data = 16'b1101010010010100;
				18'b010100110010011000: oled_data = 16'b1101010010010101;
				18'b010100110100011000: oled_data = 16'b1101110011010101;
				18'b010100110110011000: oled_data = 16'b1101110011010101;
				18'b010100111000011000: oled_data = 16'b1101110011010101;
				18'b010100111010011000: oled_data = 16'b1101110011010101;
				18'b010100111100011000: oled_data = 16'b1101110011010101;
				18'b010100111110011000: oled_data = 16'b1101110011010110;
				18'b010101000000011000: oled_data = 16'b1101010001110100;
				18'b010101000010011000: oled_data = 16'b1101110010110101;
				18'b010101000100011000: oled_data = 16'b1101110011010101;
				18'b010101000110011000: oled_data = 16'b1101110011010101;
				18'b010101001000011000: oled_data = 16'b1101110011010110;
				18'b010101001010011000: oled_data = 16'b1101010011010100;
				18'b010101001100011000: oled_data = 16'b1101010101010101;
				18'b010101001110011000: oled_data = 16'b1101110011010101;
				18'b010101010000011000: oled_data = 16'b1101110011010101;
				18'b010101010010011000: oled_data = 16'b1101110011010101;
				18'b010101010100011000: oled_data = 16'b1101010100010110;
				18'b010101010110011000: oled_data = 16'b1101110011110110;
				18'b010101011000011000: oled_data = 16'b1101110011010110;
				18'b010101011010011000: oled_data = 16'b1101110011010101;
				18'b010101011100011000: oled_data = 16'b1110010011010101;
				18'b010101011110011000: oled_data = 16'b1101110011010101;
				18'b010101100000011000: oled_data = 16'b1110010011010110;
				18'b010101100010011000: oled_data = 16'b1110010011010110;
				18'b010101100100011000: oled_data = 16'b1110010011010110;
				18'b010101100110011000: oled_data = 16'b1101110011010110;
				18'b010101101000011000: oled_data = 16'b1101010010010100;
				18'b010101101010011000: oled_data = 16'b1100110010010100;
				18'b010101101100011000: oled_data = 16'b1100010001110011;
				18'b010101101110011000: oled_data = 16'b1110010100010110;
				18'b010101110000011000: oled_data = 16'b1101110011010101;
				18'b010101110010011000: oled_data = 16'b0101100110101000;
				18'b010101110100011000: oled_data = 16'b1010110011110011;
				18'b010101110110011000: oled_data = 16'b1101110101010111;
				18'b010101111000011000: oled_data = 16'b1101110010110110;
				18'b010101111010011000: oled_data = 16'b1101110011010101;
				18'b010101111100011000: oled_data = 16'b1011101110110001;
				18'b010101111110011000: oled_data = 16'b1011001101110001;
				18'b010110000000011000: oled_data = 16'b1100110001010011;
				18'b010110000010011000: oled_data = 16'b1101110010110101;
				18'b010110000100011000: oled_data = 16'b1101010010010011;
				18'b010110000110011000: oled_data = 16'b1110110100010100;
				18'b010110001000011000: oled_data = 16'b1100101101101101;
				18'b010110001010011000: oled_data = 16'b1011001000101001;
				18'b010110001100011000: oled_data = 16'b1011101001001001;
				18'b010110001110011000: oled_data = 16'b1011001001001001;
				18'b010110010000011000: oled_data = 16'b1011001001001001;
				18'b010110010010011000: oled_data = 16'b1011001001001001;
				18'b010110010100011000: oled_data = 16'b1011001001001001;
				18'b010110010110011000: oled_data = 16'b1011001000101001;
				18'b010110011000011000: oled_data = 16'b1010101000001000;
				18'b010110011010011000: oled_data = 16'b1011001000101001;
				18'b010110011100011000: oled_data = 16'b1011001001001001;
				18'b010110011110011000: oled_data = 16'b1011001000101001;
				18'b010110100000011000: oled_data = 16'b1011001000101001;
				18'b010110100010011000: oled_data = 16'b1011001000101001;
				18'b010110100100011000: oled_data = 16'b1011001000101000;
				18'b010110100110011000: oled_data = 16'b1010101000001000;
				18'b010100011000011001: oled_data = 16'b1100010111001110;
				18'b010100011010011001: oled_data = 16'b1100110110101101;
				18'b010100011100011001: oled_data = 16'b1011010100001001;
				18'b010100011110011001: oled_data = 16'b1010110010100111;
				18'b010100100000011001: oled_data = 16'b1011110101001001;
				18'b010100100010011001: oled_data = 16'b1101010111101011;
				18'b010100100100011001: oled_data = 16'b1100110001110000;
				18'b010100100110011001: oled_data = 16'b1101110010010101;
				18'b010100101000011001: oled_data = 16'b1101010010010101;
				18'b010100101010011001: oled_data = 16'b1101110011010110;
				18'b010100101100011001: oled_data = 16'b1101110011010110;
				18'b010100101110011001: oled_data = 16'b1101010001110100;
				18'b010100110000011001: oled_data = 16'b1101110011010101;
				18'b010100110010011001: oled_data = 16'b1101010010010100;
				18'b010100110100011001: oled_data = 16'b1101110011010101;
				18'b010100110110011001: oled_data = 16'b1101110011010101;
				18'b010100111000011001: oled_data = 16'b1101110011010101;
				18'b010100111010011001: oled_data = 16'b1101110011010101;
				18'b010100111100011001: oled_data = 16'b1101110011010101;
				18'b010100111110011001: oled_data = 16'b1101110011010101;
				18'b010101000000011001: oled_data = 16'b1101010001110100;
				18'b010101000010011001: oled_data = 16'b1101110011010101;
				18'b010101000100011001: oled_data = 16'b1101110011010101;
				18'b010101000110011001: oled_data = 16'b1101110011010101;
				18'b010101001000011001: oled_data = 16'b1101110010110101;
				18'b010101001010011001: oled_data = 16'b1100110100010100;
				18'b010101001100011001: oled_data = 16'b1101111000111000;
				18'b010101001110011001: oled_data = 16'b1101110010110101;
				18'b010101010000011001: oled_data = 16'b1101110011010110;
				18'b010101010010011001: oled_data = 16'b1101110010110101;
				18'b010101010100011001: oled_data = 16'b1101110111011000;
				18'b010101010110011001: oled_data = 16'b1101110011110110;
				18'b010101011000011001: oled_data = 16'b1101110011010101;
				18'b010101011010011001: oled_data = 16'b1101110011010101;
				18'b010101011100011001: oled_data = 16'b1101110011010101;
				18'b010101011110011001: oled_data = 16'b1101110011010101;
				18'b010101100000011001: oled_data = 16'b1101110011010101;
				18'b010101100010011001: oled_data = 16'b1101110011010101;
				18'b010101100100011001: oled_data = 16'b1101110011010101;
				18'b010101100110011001: oled_data = 16'b1101110011010101;
				18'b010101101000011001: oled_data = 16'b1101010010110101;
				18'b010101101010011001: oled_data = 16'b1101010011010101;
				18'b010101101100011001: oled_data = 16'b1101010101010110;
				18'b010101101110011001: oled_data = 16'b1110010100110110;
				18'b010101110000011001: oled_data = 16'b1010101111010001;
				18'b010101110010011001: oled_data = 16'b0101000111101000;
				18'b010101110100011001: oled_data = 16'b1101011001011001;
				18'b010101110110011001: oled_data = 16'b1101010100110110;
				18'b010101111000011001: oled_data = 16'b1110010011010110;
				18'b010101111010011001: oled_data = 16'b1101010001110100;
				18'b010101111100011001: oled_data = 16'b1011001101110001;
				18'b010101111110011001: oled_data = 16'b1011001101110001;
				18'b010110000000011001: oled_data = 16'b1100110001010100;
				18'b010110000010011001: oled_data = 16'b1101010001110011;
				18'b010110000100011001: oled_data = 16'b1110010011110100;
				18'b010110000110011001: oled_data = 16'b1101110001110010;
				18'b010110001000011001: oled_data = 16'b1011101001101010;
				18'b010110001010011001: oled_data = 16'b1011001001001001;
				18'b010110001100011001: oled_data = 16'b1011001001001001;
				18'b010110001110011001: oled_data = 16'b1011001001001001;
				18'b010110010000011001: oled_data = 16'b1011001001001001;
				18'b010110010010011001: oled_data = 16'b1011001001001001;
				18'b010110010100011001: oled_data = 16'b1011001000101001;
				18'b010110010110011001: oled_data = 16'b1010101000001000;
				18'b010110011000011001: oled_data = 16'b1011001000101001;
				18'b010110011010011001: oled_data = 16'b1011001001001001;
				18'b010110011100011001: oled_data = 16'b1011001000101001;
				18'b010110011110011001: oled_data = 16'b1011001000101001;
				18'b010110100000011001: oled_data = 16'b1011001000101001;
				18'b010110100010011001: oled_data = 16'b1011001000101000;
				18'b010110100100011001: oled_data = 16'b1011001000101000;
				18'b010110100110011001: oled_data = 16'b1010101000101000;
				18'b010100011000011010: oled_data = 16'b1010010010100111;
				18'b010100011010011010: oled_data = 16'b1010010010100111;
				18'b010100011100011010: oled_data = 16'b1010110010100111;
				18'b010100011110011010: oled_data = 16'b1010110010101000;
				18'b010100100000011010: oled_data = 16'b1010110011001000;
				18'b010100100010011010: oled_data = 16'b1100110111101011;
				18'b010100100100011010: oled_data = 16'b1101010011110010;
				18'b010100100110011010: oled_data = 16'b1101010001110101;
				18'b010100101000011010: oled_data = 16'b1101110011010101;
				18'b010100101010011010: oled_data = 16'b1101110011010101;
				18'b010100101100011010: oled_data = 16'b1101110011010101;
				18'b010100101110011010: oled_data = 16'b1101010010010101;
				18'b010100110000011010: oled_data = 16'b1101110011010110;
				18'b010100110010011010: oled_data = 16'b1101110010010101;
				18'b010100110100011010: oled_data = 16'b1101110011010101;
				18'b010100110110011010: oled_data = 16'b1101110011010101;
				18'b010100111000011010: oled_data = 16'b1101110011010101;
				18'b010100111010011010: oled_data = 16'b1101110011010101;
				18'b010100111100011010: oled_data = 16'b1101110011010101;
				18'b010100111110011010: oled_data = 16'b1101110011010101;
				18'b010101000000011010: oled_data = 16'b1101010010010100;
				18'b010101000010011010: oled_data = 16'b1101110011010101;
				18'b010101000100011010: oled_data = 16'b1101110011010101;
				18'b010101000110011010: oled_data = 16'b1101110011010101;
				18'b010101001000011010: oled_data = 16'b1101110010010101;
				18'b010101001010011010: oled_data = 16'b1101110111111000;
				18'b010101001100011010: oled_data = 16'b1110011001111001;
				18'b010101001110011010: oled_data = 16'b1101110010110101;
				18'b010101010000011010: oled_data = 16'b1110010011010110;
				18'b010101010010011010: oled_data = 16'b1101010011010101;
				18'b010101010100011010: oled_data = 16'b1110011001011001;
				18'b010101010110011010: oled_data = 16'b1101110011110110;
				18'b010101011000011010: oled_data = 16'b1110010011010110;
				18'b010101011010011010: oled_data = 16'b1101110011010101;
				18'b010101011100011010: oled_data = 16'b1101110010110101;
				18'b010101011110011010: oled_data = 16'b1101110011010101;
				18'b010101100000011010: oled_data = 16'b1101110011010101;
				18'b010101100010011010: oled_data = 16'b1101110011010101;
				18'b010101100100011010: oled_data = 16'b1101110011010101;
				18'b010101100110011010: oled_data = 16'b1101110010110101;
				18'b010101101000011010: oled_data = 16'b1101110011010101;
				18'b010101101010011010: oled_data = 16'b1101110100010110;
				18'b010101101100011010: oled_data = 16'b1101110101010111;
				18'b010101101110011010: oled_data = 16'b1101110100010110;
				18'b010101110000011010: oled_data = 16'b0111101001001011;
				18'b010101110010011010: oled_data = 16'b0111101101001101;
				18'b010101110100011010: oled_data = 16'b1110011100011011;
				18'b010101110110011010: oled_data = 16'b1101010100010110;
				18'b010101111000011010: oled_data = 16'b1110010011010110;
				18'b010101111010011010: oled_data = 16'b1100110000010011;
				18'b010101111100011010: oled_data = 16'b1011001101110001;
				18'b010101111110011010: oled_data = 16'b1011001101110001;
				18'b010110000000011010: oled_data = 16'b1100010000010010;
				18'b010110000010011010: oled_data = 16'b1101110010110011;
				18'b010110000100011010: oled_data = 16'b1110110100010100;
				18'b010110000110011010: oled_data = 16'b1100101100101101;
				18'b010110001000011010: oled_data = 16'b1011001001001001;
				18'b010110001010011010: oled_data = 16'b1011001001001001;
				18'b010110001100011010: oled_data = 16'b1011001001001001;
				18'b010110001110011010: oled_data = 16'b1011001001001001;
				18'b010110010000011010: oled_data = 16'b1011001001001001;
				18'b010110010010011010: oled_data = 16'b1011001001001001;
				18'b010110010100011010: oled_data = 16'b1010101000001000;
				18'b010110010110011010: oled_data = 16'b1011001000101001;
				18'b010110011000011010: oled_data = 16'b1011001001001001;
				18'b010110011010011010: oled_data = 16'b1011001001001001;
				18'b010110011100011010: oled_data = 16'b1011001000101001;
				18'b010110011110011010: oled_data = 16'b1011001000101001;
				18'b010110100000011010: oled_data = 16'b1011001000101001;
				18'b010110100010011010: oled_data = 16'b1011001000101000;
				18'b010110100100011010: oled_data = 16'b1011001000101000;
				18'b010110100110011010: oled_data = 16'b1010101000101000;
				18'b010100011000011011: oled_data = 16'b1010110010100111;
				18'b010100011010011011: oled_data = 16'b1010110010100111;
				18'b010100011100011011: oled_data = 16'b1010110010100111;
				18'b010100011110011011: oled_data = 16'b1010110010100111;
				18'b010100100000011011: oled_data = 16'b1010110010100111;
				18'b010100100010011011: oled_data = 16'b1100110110001011;
				18'b010100100100011011: oled_data = 16'b1101010011110011;
				18'b010100100110011011: oled_data = 16'b1101010001110101;
				18'b010100101000011011: oled_data = 16'b1110010011010110;
				18'b010100101010011011: oled_data = 16'b1101110011010101;
				18'b010100101100011011: oled_data = 16'b1101010010010100;
				18'b010100101110011011: oled_data = 16'b1101110010110101;
				18'b010100110000011011: oled_data = 16'b1101110011010101;
				18'b010100110010011011: oled_data = 16'b1101110010010101;
				18'b010100110100011011: oled_data = 16'b1101110011010110;
				18'b010100110110011011: oled_data = 16'b1110010011010110;
				18'b010100111000011011: oled_data = 16'b1101110011010101;
				18'b010100111010011011: oled_data = 16'b1101110011010101;
				18'b010100111100011011: oled_data = 16'b1110010011010110;
				18'b010100111110011011: oled_data = 16'b1101110010110101;
				18'b010101000000011011: oled_data = 16'b1101010010010100;
				18'b010101000010011011: oled_data = 16'b1101110011010110;
				18'b010101000100011011: oled_data = 16'b1101110011010101;
				18'b010101000110011011: oled_data = 16'b1101110011010101;
				18'b010101001000011011: oled_data = 16'b1101010011010100;
				18'b010101001010011011: oled_data = 16'b1110011010111010;
				18'b010101001100011011: oled_data = 16'b1101111001111000;
				18'b010101001110011011: oled_data = 16'b1101010011010101;
				18'b010101010000011011: oled_data = 16'b1101110011010101;
				18'b010101010010011011: oled_data = 16'b1101110100010110;
				18'b010101010100011011: oled_data = 16'b1110011001011001;
				18'b010101010110011011: oled_data = 16'b1101110011010101;
				18'b010101011000011011: oled_data = 16'b1110010011110110;
				18'b010101011010011011: oled_data = 16'b1101010001110100;
				18'b010101011100011011: oled_data = 16'b1101110010110101;
				18'b010101011110011011: oled_data = 16'b1101110011010101;
				18'b010101100000011011: oled_data = 16'b1101110011010101;
				18'b010101100010011011: oled_data = 16'b1101110011010101;
				18'b010101100100011011: oled_data = 16'b1101110011010110;
				18'b010101100110011011: oled_data = 16'b1101010001110100;
				18'b010101101000011011: oled_data = 16'b1101010011010101;
				18'b010101101010011011: oled_data = 16'b1101110110010111;
				18'b010101101100011011: oled_data = 16'b1101110100110110;
				18'b010101101110011011: oled_data = 16'b1100110010010100;
				18'b010101110000011011: oled_data = 16'b0101100111001000;
				18'b010101110010011011: oled_data = 16'b1011010101010100;
				18'b010101110100011011: oled_data = 16'b1110011011111010;
				18'b010101110110011011: oled_data = 16'b1100110011110101;
				18'b010101111000011011: oled_data = 16'b1101010011110101;
				18'b010101111010011011: oled_data = 16'b1101110111111000;
				18'b010101111100011011: oled_data = 16'b1011001111110010;
				18'b010101111110011011: oled_data = 16'b1011001101110001;
				18'b010110000000011011: oled_data = 16'b1011101111010001;
				18'b010110000010011011: oled_data = 16'b1110110100010100;
				18'b010110000100011011: oled_data = 16'b1101110001110001;
				18'b010110000110011011: oled_data = 16'b1011101001101010;
				18'b010110001000011011: oled_data = 16'b1011101001001001;
				18'b010110001010011011: oled_data = 16'b1100001011001100;
				18'b010110001100011011: oled_data = 16'b1011101001101010;
				18'b010110001110011011: oled_data = 16'b1011001001001001;
				18'b010110010000011011: oled_data = 16'b1011001001001001;
				18'b010110010010011011: oled_data = 16'b1011001000101000;
				18'b010110010100011011: oled_data = 16'b1010101000101001;
				18'b010110010110011011: oled_data = 16'b1011001001001001;
				18'b010110011000011011: oled_data = 16'b1011001001001001;
				18'b010110011010011011: oled_data = 16'b1011001000101001;
				18'b010110011100011011: oled_data = 16'b1011001000101001;
				18'b010110011110011011: oled_data = 16'b1011001000101001;
				18'b010110100000011011: oled_data = 16'b1011001000101001;
				18'b010110100010011011: oled_data = 16'b1011001000101000;
				18'b010110100100011011: oled_data = 16'b1011001000101000;
				18'b010110100110011011: oled_data = 16'b1010101000101000;
				18'b010100011000011100: oled_data = 16'b1010110010100111;
				18'b010100011010011100: oled_data = 16'b1010110010100111;
				18'b010100011100011100: oled_data = 16'b1010110010100111;
				18'b010100011110011100: oled_data = 16'b1010110010100111;
				18'b010100100000011100: oled_data = 16'b1010110010100111;
				18'b010100100010011100: oled_data = 16'b1100110110001010;
				18'b010100100100011100: oled_data = 16'b1101010011110011;
				18'b010100100110011100: oled_data = 16'b1101010010010101;
				18'b010100101000011100: oled_data = 16'b1101110011010110;
				18'b010100101010011100: oled_data = 16'b1101110011010101;
				18'b010100101100011100: oled_data = 16'b1101010010010100;
				18'b010100101110011100: oled_data = 16'b1101110011110110;
				18'b010100110000011100: oled_data = 16'b1101110011010101;
				18'b010100110010011100: oled_data = 16'b1101010010010101;
				18'b010100110100011100: oled_data = 16'b1110010011010110;
				18'b010100110110011100: oled_data = 16'b1110010011010110;
				18'b010100111000011100: oled_data = 16'b1101110011010101;
				18'b010100111010011100: oled_data = 16'b1101110011010101;
				18'b010100111100011100: oled_data = 16'b1110010011110110;
				18'b010100111110011100: oled_data = 16'b1101110010110101;
				18'b010101000000011100: oled_data = 16'b1101110010010101;
				18'b010101000010011100: oled_data = 16'b1101110011010110;
				18'b010101000100011100: oled_data = 16'b1101110011010101;
				18'b010101000110011100: oled_data = 16'b1101110010110101;
				18'b010101001000011100: oled_data = 16'b1101110101110110;
				18'b010101001010011100: oled_data = 16'b1110111100011011;
				18'b010101001100011100: oled_data = 16'b1101011001111000;
				18'b010101001110011100: oled_data = 16'b1101010011010101;
				18'b010101010000011100: oled_data = 16'b1101110010110101;
				18'b010101010010011100: oled_data = 16'b1101110110010111;
				18'b010101010100011100: oled_data = 16'b1110011010111010;
				18'b010101010110011100: oled_data = 16'b1101110011010101;
				18'b010101011000011100: oled_data = 16'b1101110010110101;
				18'b010101011010011100: oled_data = 16'b1101010010010100;
				18'b010101011100011100: oled_data = 16'b1101110011010101;
				18'b010101011110011100: oled_data = 16'b1101110011010101;
				18'b010101100000011100: oled_data = 16'b1101110011010101;
				18'b010101100010011100: oled_data = 16'b1101110011010101;
				18'b010101100100011100: oled_data = 16'b1101110010110101;
				18'b010101100110011100: oled_data = 16'b1101010001110100;
				18'b010101101000011100: oled_data = 16'b1101110011110110;
				18'b010101101010011100: oled_data = 16'b1101110111111001;
				18'b010101101100011100: oled_data = 16'b1101110100110110;
				18'b010101101110011100: oled_data = 16'b1001101101001111;
				18'b010101110000011100: oled_data = 16'b0101001001001001;
				18'b010101110010011100: oled_data = 16'b1101111011011001;
				18'b010101110100011100: oled_data = 16'b1101111010111001;
				18'b010101110110011100: oled_data = 16'b1100110010110101;
				18'b010101111000011100: oled_data = 16'b1101010110010111;
				18'b010101111010011100: oled_data = 16'b1110111100011011;
				18'b010101111100011100: oled_data = 16'b1100010011110100;
				18'b010101111110011100: oled_data = 16'b1010101100110000;
				18'b010110000000011100: oled_data = 16'b1100110000110001;
				18'b010110000010011100: oled_data = 16'b1110110100010100;
				18'b010110000100011100: oled_data = 16'b1100101101101101;
				18'b010110000110011100: oled_data = 16'b1011001000101001;
				18'b010110001000011100: oled_data = 16'b1011101010001010;
				18'b010110001010011100: oled_data = 16'b1101001110001110;
				18'b010110001100011100: oled_data = 16'b1011001001001010;
				18'b010110001110011100: oled_data = 16'b1011101001001001;
				18'b010110010000011100: oled_data = 16'b1011001001001001;
				18'b010110010010011100: oled_data = 16'b1010101000001000;
				18'b010110010100011100: oled_data = 16'b1011101001001001;
				18'b010110010110011100: oled_data = 16'b1011001001001001;
				18'b010110011000011100: oled_data = 16'b1010000111101000;
				18'b010110011010011100: oled_data = 16'b1010000111000111;
				18'b010110011100011100: oled_data = 16'b1011001001001001;
				18'b010110011110011100: oled_data = 16'b1011001000101000;
				18'b010110100000011100: oled_data = 16'b1011001000101001;
				18'b010110100010011100: oled_data = 16'b1011001000101000;
				18'b010110100100011100: oled_data = 16'b1011001000101000;
				18'b010110100110011100: oled_data = 16'b1010101000101000;
				18'b010100011000011101: oled_data = 16'b1010110010100111;
				18'b010100011010011101: oled_data = 16'b1010110010100111;
				18'b010100011100011101: oled_data = 16'b1010110010100111;
				18'b010100011110011101: oled_data = 16'b1010110010100111;
				18'b010100100000011101: oled_data = 16'b1010110010100111;
				18'b010100100010011101: oled_data = 16'b1100010110001010;
				18'b010100100100011101: oled_data = 16'b1101010011010011;
				18'b010100100110011101: oled_data = 16'b1101110010110101;
				18'b010100101000011101: oled_data = 16'b1101110011010110;
				18'b010100101010011101: oled_data = 16'b1101110010010101;
				18'b010100101100011101: oled_data = 16'b1101010010010100;
				18'b010100101110011101: oled_data = 16'b1101110011010110;
				18'b010100110000011101: oled_data = 16'b1101110011010101;
				18'b010100110010011101: oled_data = 16'b1101010001010100;
				18'b010100110100011101: oled_data = 16'b1101110011010101;
				18'b010100110110011101: oled_data = 16'b1101110011010110;
				18'b010100111000011101: oled_data = 16'b1101110011010101;
				18'b010100111010011101: oled_data = 16'b1101110011010101;
				18'b010100111100011101: oled_data = 16'b1101110011010101;
				18'b010100111110011101: oled_data = 16'b1101010010010100;
				18'b010101000000011101: oled_data = 16'b1101110010110101;
				18'b010101000010011101: oled_data = 16'b1101110011010110;
				18'b010101000100011101: oled_data = 16'b1101110011010101;
				18'b010101000110011101: oled_data = 16'b1101010011010101;
				18'b010101001000011101: oled_data = 16'b1110011010011001;
				18'b010101001010011101: oled_data = 16'b1110111100111011;
				18'b010101001100011101: oled_data = 16'b1101111001011000;
				18'b010101001110011101: oled_data = 16'b1101010011010101;
				18'b010101010000011101: oled_data = 16'b1101110011010101;
				18'b010101010010011101: oled_data = 16'b1101111000111000;
				18'b010101010100011101: oled_data = 16'b1110011010111010;
				18'b010101010110011101: oled_data = 16'b1101010010110101;
				18'b010101011000011101: oled_data = 16'b1101010001110100;
				18'b010101011010011101: oled_data = 16'b1101110010110101;
				18'b010101011100011101: oled_data = 16'b1101110011010101;
				18'b010101011110011101: oled_data = 16'b1101110011010101;
				18'b010101100000011101: oled_data = 16'b1101110010110101;
				18'b010101100010011101: oled_data = 16'b1101110011010101;
				18'b010101100100011101: oled_data = 16'b1101010010010100;
				18'b010101100110011101: oled_data = 16'b1101110010010101;
				18'b010101101000011101: oled_data = 16'b1101110100110110;
				18'b010101101010011101: oled_data = 16'b1110011000011001;
				18'b010101101100011101: oled_data = 16'b1101010011110101;
				18'b010101101110011101: oled_data = 16'b0110101001001010;
				18'b010101110000011101: oled_data = 16'b1000101111110000;
				18'b010101110010011101: oled_data = 16'b1111011101011011;
				18'b010101110100011101: oled_data = 16'b1101111000111000;
				18'b010101110110011101: oled_data = 16'b1101010101110110;
				18'b010101111000011101: oled_data = 16'b1110111011011011;
				18'b010101111010011101: oled_data = 16'b1110111100011011;
				18'b010101111100011101: oled_data = 16'b1101111000111001;
				18'b010101111110011101: oled_data = 16'b1011001110010000;
				18'b010110000000011101: oled_data = 16'b1110010011010100;
				18'b010110000010011101: oled_data = 16'b1110010011010011;
				18'b010110000100011101: oled_data = 16'b1011101010001010;
				18'b010110000110011101: oled_data = 16'b1011001000101001;
				18'b010110001000011101: oled_data = 16'b1100001011101011;
				18'b010110001010011101: oled_data = 16'b1100001100101100;
				18'b010110001100011101: oled_data = 16'b1011001000101001;
				18'b010110001110011101: oled_data = 16'b1011101001001001;
				18'b010110010000011101: oled_data = 16'b1011001000101000;
				18'b010110010010011101: oled_data = 16'b1011001001001001;
				18'b010110010100011101: oled_data = 16'b1011101001001001;
				18'b010110010110011101: oled_data = 16'b1010001000001000;
				18'b010110011000011101: oled_data = 16'b1001000101100110;
				18'b010110011010011101: oled_data = 16'b1010101000001000;
				18'b010110011100011101: oled_data = 16'b1011001000101001;
				18'b010110011110011101: oled_data = 16'b1011001000101000;
				18'b010110100000011101: oled_data = 16'b1011001000101001;
				18'b010110100010011101: oled_data = 16'b1011001000101000;
				18'b010110100100011101: oled_data = 16'b1011001000101000;
				18'b010110100110011101: oled_data = 16'b1010101000101000;
				18'b010100011000011110: oled_data = 16'b1010110010100111;
				18'b010100011010011110: oled_data = 16'b1010110010100111;
				18'b010100011100011110: oled_data = 16'b1010110010100111;
				18'b010100011110011110: oled_data = 16'b1010110010100111;
				18'b010100100000011110: oled_data = 16'b1010110011000111;
				18'b010100100010011110: oled_data = 16'b1100110110001101;
				18'b010100100100011110: oled_data = 16'b1100110010010011;
				18'b010100100110011110: oled_data = 16'b1110010011010101;
				18'b010100101000011110: oled_data = 16'b1110010011010110;
				18'b010100101010011110: oled_data = 16'b1101010001110100;
				18'b010100101100011110: oled_data = 16'b1101110010110101;
				18'b010100101110011110: oled_data = 16'b1101110011010101;
				18'b010100110000011110: oled_data = 16'b1101110011010101;
				18'b010100110010011110: oled_data = 16'b1101010010010100;
				18'b010100110100011110: oled_data = 16'b1101110010110101;
				18'b010100110110011110: oled_data = 16'b1101110011010110;
				18'b010100111000011110: oled_data = 16'b1101110011010101;
				18'b010100111010011110: oled_data = 16'b1101110011010110;
				18'b010100111100011110: oled_data = 16'b1101110010010101;
				18'b010100111110011110: oled_data = 16'b1101010010010100;
				18'b010101000000011110: oled_data = 16'b1101110010110101;
				18'b010101000010011110: oled_data = 16'b1101110011010101;
				18'b010101000100011110: oled_data = 16'b1101110011010101;
				18'b010101000110011110: oled_data = 16'b1101010100010101;
				18'b010101001000011110: oled_data = 16'b1111011100011011;
				18'b010101001010011110: oled_data = 16'b1110111100011011;
				18'b010101001100011110: oled_data = 16'b1110011010011001;
				18'b010101001110011110: oled_data = 16'b1101010011110101;
				18'b010101010000011110: oled_data = 16'b1101110011010101;
				18'b010101010010011110: oled_data = 16'b1110011010011010;
				18'b010101010100011110: oled_data = 16'b1101111001111001;
				18'b010101010110011110: oled_data = 16'b1100110001010011;
				18'b010101011000011110: oled_data = 16'b1101110010110101;
				18'b010101011010011110: oled_data = 16'b1101110011010110;
				18'b010101011100011110: oled_data = 16'b1101110011010101;
				18'b010101011110011110: oled_data = 16'b1101110011010101;
				18'b010101100000011110: oled_data = 16'b1101110010110101;
				18'b010101100010011110: oled_data = 16'b1101110011010101;
				18'b010101100100011110: oled_data = 16'b1101010010010100;
				18'b010101100110011110: oled_data = 16'b1101110010110101;
				18'b010101101000011110: oled_data = 16'b1110010110111000;
				18'b010101101010011110: oled_data = 16'b1101010110110111;
				18'b010101101100011110: oled_data = 16'b1011110100010101;
				18'b010101101110011110: oled_data = 16'b0101101001001001;
				18'b010101110000011110: oled_data = 16'b1101011000011000;
				18'b010101110010011110: oled_data = 16'b1110111100011011;
				18'b010101110100011110: oled_data = 16'b1100110111110110;
				18'b010101110110011110: oled_data = 16'b1101011001111000;
				18'b010101111000011110: oled_data = 16'b1100111000111000;
				18'b010101111010011110: oled_data = 16'b1101011010011001;
				18'b010101111100011110: oled_data = 16'b1101111010011010;
				18'b010101111110011110: oled_data = 16'b1100110010010011;
				18'b010110000000011110: oled_data = 16'b1110110100010100;
				18'b010110000010011110: oled_data = 16'b1101001111110000;
				18'b010110000100011110: oled_data = 16'b1011001000101001;
				18'b010110000110011110: oled_data = 16'b1011101001001001;
				18'b010110001000011110: oled_data = 16'b1100001100001100;
				18'b010110001010011110: oled_data = 16'b1011101010001010;
				18'b010110001100011110: oled_data = 16'b1011001001001001;
				18'b010110001110011110: oled_data = 16'b1011001001001001;
				18'b010110010000011110: oled_data = 16'b1010101000101000;
				18'b010110010010011110: oled_data = 16'b1011001001001001;
				18'b010110010100011110: oled_data = 16'b1010101000101000;
				18'b010110010110011110: oled_data = 16'b1000100101100110;
				18'b010110011000011110: oled_data = 16'b1001100110100111;
				18'b010110011010011110: oled_data = 16'b1011101010001010;
				18'b010110011100011110: oled_data = 16'b1011101010101010;
				18'b010110011110011110: oled_data = 16'b1011001000101000;
				18'b010110100000011110: oled_data = 16'b1011001000101001;
				18'b010110100010011110: oled_data = 16'b1011001000101000;
				18'b010110100100011110: oled_data = 16'b1011001000101000;
				18'b010110100110011110: oled_data = 16'b1010101000101000;
				18'b010100011000011111: oled_data = 16'b1011110101001001;
				18'b010100011010011111: oled_data = 16'b1011010100101000;
				18'b010100011100011111: oled_data = 16'b1011010011100111;
				18'b010100011110011111: oled_data = 16'b1010110011100111;
				18'b010100100000011111: oled_data = 16'b1100010110001001;
				18'b010100100010011111: oled_data = 16'b1101010110010000;
				18'b010100100100011111: oled_data = 16'b1101010010010100;
				18'b010100100110011111: oled_data = 16'b1101110011010101;
				18'b010100101000011111: oled_data = 16'b1101110010110101;
				18'b010100101010011111: oled_data = 16'b1101010001110100;
				18'b010100101100011111: oled_data = 16'b1101110011010101;
				18'b010100101110011111: oled_data = 16'b1110010011010101;
				18'b010100110000011111: oled_data = 16'b1110010011010110;
				18'b010100110010011111: oled_data = 16'b1101110010010101;
				18'b010100110100011111: oled_data = 16'b1101110010010101;
				18'b010100110110011111: oled_data = 16'b1110010011010110;
				18'b010100111000011111: oled_data = 16'b1101110011010101;
				18'b010100111010011111: oled_data = 16'b1101110011010101;
				18'b010100111100011111: oled_data = 16'b1101010010010100;
				18'b010100111110011111: oled_data = 16'b1100110010010100;
				18'b010101000000011111: oled_data = 16'b1101110011010101;
				18'b010101000010011111: oled_data = 16'b1101110011010110;
				18'b010101000100011111: oled_data = 16'b1101110010110101;
				18'b010101000110011111: oled_data = 16'b1110010111111000;
				18'b010101001000011111: oled_data = 16'b1110111100011011;
				18'b010101001010011111: oled_data = 16'b1110111100011011;
				18'b010101001100011111: oled_data = 16'b1110011010111010;
				18'b010101001110011111: oled_data = 16'b1101010011110101;
				18'b010101010000011111: oled_data = 16'b1101010100010110;
				18'b010101010010011111: oled_data = 16'b1110011010111010;
				18'b010101010100011111: oled_data = 16'b1101011000011000;
				18'b010101010110011111: oled_data = 16'b1101010010110101;
				18'b010101011000011111: oled_data = 16'b1101110011010110;
				18'b010101011010011111: oled_data = 16'b1101110011010101;
				18'b010101011100011111: oled_data = 16'b1101110011010101;
				18'b010101011110011111: oled_data = 16'b1101110011010101;
				18'b010101100000011111: oled_data = 16'b1101110011010101;
				18'b010101100010011111: oled_data = 16'b1101110010110101;
				18'b010101100100011111: oled_data = 16'b1101010010010101;
				18'b010101100110011111: oled_data = 16'b1101010011110101;
				18'b010101101000011111: oled_data = 16'b1110011010011010;
				18'b010101101010011111: oled_data = 16'b1101011000111000;
				18'b010101101100011111: oled_data = 16'b1011010100010100;
				18'b010101101110011111: oled_data = 16'b0100000110000110;
				18'b010101110000011111: oled_data = 16'b0110001010101011;
				18'b010101110010011111: oled_data = 16'b0101101001101001;
				18'b010101110100011111: oled_data = 16'b0101001000101000;
				18'b010101110110011111: oled_data = 16'b0100101000000111;
				18'b010101111000011111: oled_data = 16'b0011100110000101;
				18'b010101111010011111: oled_data = 16'b0100000111100111;
				18'b010101111100011111: oled_data = 16'b0110001001101010;
				18'b010101111110011111: oled_data = 16'b1100110010110011;
				18'b010110000000011111: oled_data = 16'b1110110100010100;
				18'b010110000010011111: oled_data = 16'b1100001100001101;
				18'b010110000100011111: oled_data = 16'b1011001000101001;
				18'b010110000110011111: oled_data = 16'b1011101001001001;
				18'b010110001000011111: oled_data = 16'b1011101010001010;
				18'b010110001010011111: oled_data = 16'b1011001001001001;
				18'b010110001100011111: oled_data = 16'b1011001001001001;
				18'b010110001110011111: oled_data = 16'b1010101000101000;
				18'b010110010000011111: oled_data = 16'b1011001001001001;
				18'b010110010010011111: oled_data = 16'b1011001000101001;
				18'b010110010100011111: oled_data = 16'b1001000110000111;
				18'b010110010110011111: oled_data = 16'b1001000101100110;
				18'b010110011000011111: oled_data = 16'b1011001001001010;
				18'b010110011010011111: oled_data = 16'b1101001111101111;
				18'b010110011100011111: oled_data = 16'b1011101010001010;
				18'b010110011110011111: oled_data = 16'b1011001000101000;
				18'b010110100000011111: oled_data = 16'b1011001000101001;
				18'b010110100010011111: oled_data = 16'b1011001000101000;
				18'b010110100100011111: oled_data = 16'b1011001000101000;
				18'b010110100110011111: oled_data = 16'b1010101000101000;
				18'b010100011000100000: oled_data = 16'b1101010110001110;
				18'b010100011010100000: oled_data = 16'b1101010111001110;
				18'b010100011100100000: oled_data = 16'b1101010110101101;
				18'b010100011110100000: oled_data = 16'b1100110110101101;
				18'b010100100000100000: oled_data = 16'b1101010111001101;
				18'b010100100010100000: oled_data = 16'b1101010011110001;
				18'b010100100100100000: oled_data = 16'b1101010010010101;
				18'b010100100110100000: oled_data = 16'b1101110010010101;
				18'b010100101000100000: oled_data = 16'b1101010010010101;
				18'b010100101010100000: oled_data = 16'b1101010010010100;
				18'b010100101100100000: oled_data = 16'b1110010011010110;
				18'b010100101110100000: oled_data = 16'b1110010011010101;
				18'b010100110000100000: oled_data = 16'b1110010011010101;
				18'b010100110010100000: oled_data = 16'b1101110010110101;
				18'b010100110100100000: oled_data = 16'b1101010001110100;
				18'b010100110110100000: oled_data = 16'b1101110011010101;
				18'b010100111000100000: oled_data = 16'b1101110011010101;
				18'b010100111010100000: oled_data = 16'b1101110010110101;
				18'b010100111100100000: oled_data = 16'b1101010010010100;
				18'b010100111110100000: oled_data = 16'b1101010011110110;
				18'b010101000000100000: oled_data = 16'b1101110011010101;
				18'b010101000010100000: oled_data = 16'b1101110011010101;
				18'b010101000100100000: oled_data = 16'b1101010011110101;
				18'b010101000110100000: oled_data = 16'b1110011010111010;
				18'b010101001000100000: oled_data = 16'b1110011100011010;
				18'b010101001010100000: oled_data = 16'b1110011011011010;
				18'b010101001100100000: oled_data = 16'b1101011001011000;
				18'b010101001110100000: oled_data = 16'b1100110010110100;
				18'b010101010000100000: oled_data = 16'b1100110011110101;
				18'b010101010010100000: oled_data = 16'b1110011011011010;
				18'b010101010100100000: oled_data = 16'b1110011010011010;
				18'b010101010110100000: oled_data = 16'b1101110011110110;
				18'b010101011000100000: oled_data = 16'b1101110011010110;
				18'b010101011010100000: oled_data = 16'b1101110011010101;
				18'b010101011100100000: oled_data = 16'b1101110011010101;
				18'b010101011110100000: oled_data = 16'b1101110011010101;
				18'b010101100000100000: oled_data = 16'b1101110011010110;
				18'b010101100010100000: oled_data = 16'b1101010001110100;
				18'b010101100100100000: oled_data = 16'b1101010010010101;
				18'b010101100110100000: oled_data = 16'b1101010110110111;
				18'b010101101000100000: oled_data = 16'b1110111100011011;
				18'b010101101010100000: oled_data = 16'b1110111101011011;
				18'b010101101100100000: oled_data = 16'b1100010111110110;
				18'b010101101110100000: oled_data = 16'b0110001010001010;
				18'b010101110000100000: oled_data = 16'b0101101001101001;
				18'b010101110010100000: oled_data = 16'b0101101010001001;
				18'b010101110100100000: oled_data = 16'b0110001010001010;
				18'b010101110110100000: oled_data = 16'b0110101011101011;
				18'b010101111000100000: oled_data = 16'b0111001101001101;
				18'b010101111010100000: oled_data = 16'b0111101110101110;
				18'b010101111100100000: oled_data = 16'b1001110000010000;
				18'b010101111110100000: oled_data = 16'b1101010011010011;
				18'b010110000000100000: oled_data = 16'b1110010011110011;
				18'b010110000010100000: oled_data = 16'b1011001001101010;
				18'b010110000100100000: oled_data = 16'b1011001000101001;
				18'b010110000110100000: oled_data = 16'b1011001001001001;
				18'b010110001000100000: oled_data = 16'b1011001001001001;
				18'b010110001010100000: oled_data = 16'b1011001001001001;
				18'b010110001100100000: oled_data = 16'b1011001001001001;
				18'b010110001110100000: oled_data = 16'b1010101000101001;
				18'b010110010000100000: oled_data = 16'b1011001001001001;
				18'b010110010010100000: oled_data = 16'b1001100110100111;
				18'b010110010100100000: oled_data = 16'b1000100101000110;
				18'b010110010110100000: oled_data = 16'b1010000111001000;
				18'b010110011000100000: oled_data = 16'b1100101101001101;
				18'b010110011010100000: oled_data = 16'b1100001100001100;
				18'b010110011100100000: oled_data = 16'b1011001000101000;
				18'b010110011110100000: oled_data = 16'b1011001000101001;
				18'b010110100000100000: oled_data = 16'b1011001000101001;
				18'b010110100010100000: oled_data = 16'b1011001000101000;
				18'b010110100100100000: oled_data = 16'b1011001000101000;
				18'b010110100110100000: oled_data = 16'b1010101000101000;
				18'b010100011000100001: oled_data = 16'b1101110011010110;
				18'b010100011010100001: oled_data = 16'b1101110011010110;
				18'b010100011100100001: oled_data = 16'b1101110011110101;
				18'b010100011110100001: oled_data = 16'b1101110011010101;
				18'b010100100000100001: oled_data = 16'b1101110011010101;
				18'b010100100010100001: oled_data = 16'b1101010010110101;
				18'b010100100100100001: oled_data = 16'b1101110010010101;
				18'b010100100110100001: oled_data = 16'b1101010010010101;
				18'b010100101000100001: oled_data = 16'b1101010010010100;
				18'b010100101010100001: oled_data = 16'b1101110010110101;
				18'b010100101100100001: oled_data = 16'b1101110011010110;
				18'b010100101110100001: oled_data = 16'b1101110011010101;
				18'b010100110000100001: oled_data = 16'b1101110011010101;
				18'b010100110010100001: oled_data = 16'b1101110011010101;
				18'b010100110100100001: oled_data = 16'b1101110010010101;
				18'b010100110110100001: oled_data = 16'b1101110011010101;
				18'b010100111000100001: oled_data = 16'b1101110011010101;
				18'b010100111010100001: oled_data = 16'b1101110010110101;
				18'b010100111100100001: oled_data = 16'b1101010010010100;
				18'b010100111110100001: oled_data = 16'b1101110101110111;
				18'b010101000000100001: oled_data = 16'b1101110011010101;
				18'b010101000010100001: oled_data = 16'b1101110010110101;
				18'b010101000100100001: oled_data = 16'b1101110110010111;
				18'b010101000110100001: oled_data = 16'b1110111100011010;
				18'b010101001000100001: oled_data = 16'b1110011011111010;
				18'b010101001010100001: oled_data = 16'b1110111011111010;
				18'b010101001100100001: oled_data = 16'b1110111100011010;
				18'b010101001110100001: oled_data = 16'b1101010101010110;
				18'b010101010000100001: oled_data = 16'b1101110110110111;
				18'b010101010010100001: oled_data = 16'b1111011100111100;
				18'b010101010100100001: oled_data = 16'b1110011010011010;
				18'b010101010110100001: oled_data = 16'b1101110011010110;
				18'b010101011000100001: oled_data = 16'b1101110011010110;
				18'b010101011010100001: oled_data = 16'b1101110011010101;
				18'b010101011100100001: oled_data = 16'b1101110011010101;
				18'b010101011110100001: oled_data = 16'b1101110011010101;
				18'b010101100000100001: oled_data = 16'b1101110010110101;
				18'b010101100010100001: oled_data = 16'b1101010001010100;
				18'b010101100100100001: oled_data = 16'b1101010100010101;
				18'b010101100110100001: oled_data = 16'b1110011011011010;
				18'b010101101000100001: oled_data = 16'b1110111100011010;
				18'b010101101010100001: oled_data = 16'b1110111100011010;
				18'b010101101100100001: oled_data = 16'b1110111100011011;
				18'b010101101110100001: oled_data = 16'b1110011011011010;
				18'b010101110000100001: oled_data = 16'b1110011011011010;
				18'b010101110010100001: oled_data = 16'b1110111011011010;
				18'b010101110100100001: oled_data = 16'b1110111011011010;
				18'b010101110110100001: oled_data = 16'b1110111011111011;
				18'b010101111000100001: oled_data = 16'b1110111100011011;
				18'b010101111010100001: oled_data = 16'b1101111010111010;
				18'b010101111100100001: oled_data = 16'b1101111000010111;
				18'b010101111110100001: oled_data = 16'b1110010100010100;
				18'b010110000000100001: oled_data = 16'b1101110001110001;
				18'b010110000010100001: oled_data = 16'b1011001000101001;
				18'b010110000100100001: oled_data = 16'b1011001001001001;
				18'b010110000110100001: oled_data = 16'b1011001001001001;
				18'b010110001000100001: oled_data = 16'b1011001001001001;
				18'b010110001010100001: oled_data = 16'b1011001001001001;
				18'b010110001100100001: oled_data = 16'b1010101000101001;
				18'b010110001110100001: oled_data = 16'b1011001001001001;
				18'b010110010000100001: oled_data = 16'b1010000111101000;
				18'b010110010010100001: oled_data = 16'b1000100101000110;
				18'b010110010100100001: oled_data = 16'b1001100110000111;
				18'b010110010110100001: oled_data = 16'b1011001000101001;
				18'b010110011000100001: oled_data = 16'b1011101010001010;
				18'b010110011010100001: oled_data = 16'b1011001001001001;
				18'b010110011100100001: oled_data = 16'b1011001000101001;
				18'b010110011110100001: oled_data = 16'b1011001000101001;
				18'b010110100000100001: oled_data = 16'b1011001000101001;
				18'b010110100010100001: oled_data = 16'b1011001000101000;
				18'b010110100100100001: oled_data = 16'b1011001000101000;
				18'b010110100110100001: oled_data = 16'b1010101000101000;
				18'b010100011000100010: oled_data = 16'b1101110011110110;
				18'b010100011010100010: oled_data = 16'b1101110011010110;
				18'b010100011100100010: oled_data = 16'b1101110011110110;
				18'b010100011110100010: oled_data = 16'b1110010011010110;
				18'b010100100000100010: oled_data = 16'b1110010011010110;
				18'b010100100010100010: oled_data = 16'b1101110010110101;
				18'b010100100100100010: oled_data = 16'b1101010001110100;
				18'b010100100110100010: oled_data = 16'b1101110010110101;
				18'b010100101000100010: oled_data = 16'b1101010001010100;
				18'b010100101010100010: oled_data = 16'b1101110011010101;
				18'b010100101100100010: oled_data = 16'b1101010010010100;
				18'b010100101110100010: oled_data = 16'b1101110011010101;
				18'b010100110000100010: oled_data = 16'b1101110011010101;
				18'b010100110010100010: oled_data = 16'b1101110011010101;
				18'b010100110100100010: oled_data = 16'b1101110011010110;
				18'b010100110110100010: oled_data = 16'b1101110011010101;
				18'b010100111000100010: oled_data = 16'b1101110011010110;
				18'b010100111010100010: oled_data = 16'b1101110010010101;
				18'b010100111100100010: oled_data = 16'b1101010011010101;
				18'b010100111110100010: oled_data = 16'b1101111000011000;
				18'b010101000000100010: oled_data = 16'b1101110011010101;
				18'b010101000010100010: oled_data = 16'b1101110011110101;
				18'b010101000100100010: oled_data = 16'b1110111010011010;
				18'b010101000110100010: oled_data = 16'b1110111100011010;
				18'b010101001000100010: oled_data = 16'b1110111011111010;
				18'b010101001010100010: oled_data = 16'b1110111011111010;
				18'b010101001100100010: oled_data = 16'b1110111100011010;
				18'b010101001110100010: oled_data = 16'b1100110110010101;
				18'b010101010000100010: oled_data = 16'b1101111000111000;
				18'b010101010010100010: oled_data = 16'b1110111100111011;
				18'b010101010100100010: oled_data = 16'b1110011010011010;
				18'b010101010110100010: oled_data = 16'b1101110011010101;
				18'b010101011000100010: oled_data = 16'b1101110011010101;
				18'b010101011010100010: oled_data = 16'b1101110011010101;
				18'b010101011100100010: oled_data = 16'b1101110011010101;
				18'b010101011110100010: oled_data = 16'b1101110011010110;
				18'b010101100000100010: oled_data = 16'b1101010001110100;
				18'b010101100010100010: oled_data = 16'b1101010010110100;
				18'b010101100100100010: oled_data = 16'b1101111000110111;
				18'b010101100110100010: oled_data = 16'b1110111100111010;
				18'b010101101000100010: oled_data = 16'b1110111100011010;
				18'b010101101010100010: oled_data = 16'b1110111100011010;
				18'b010101101100100010: oled_data = 16'b1110111100011011;
				18'b010101101110100010: oled_data = 16'b1110111100011011;
				18'b010101110000100010: oled_data = 16'b1110111100011010;
				18'b010101110010100010: oled_data = 16'b1110111100011011;
				18'b010101110100100010: oled_data = 16'b1110111100011010;
				18'b010101110110100010: oled_data = 16'b1110111100011010;
				18'b010101111000100010: oled_data = 16'b1101111010111001;
				18'b010101111010100010: oled_data = 16'b1110011011011010;
				18'b010101111100100010: oled_data = 16'b1101110110110110;
				18'b010101111110100010: oled_data = 16'b1110010100010100;
				18'b010110000000100010: oled_data = 16'b1100101111001111;
				18'b010110000010100010: oled_data = 16'b1011001000001000;
				18'b010110000100100010: oled_data = 16'b1011101001001001;
				18'b010110000110100010: oled_data = 16'b1011001001001001;
				18'b010110001000100010: oled_data = 16'b1011001001001001;
				18'b010110001010100010: oled_data = 16'b1011001001001001;
				18'b010110001100100010: oled_data = 16'b1010101000101000;
				18'b010110001110100010: oled_data = 16'b1011001001001001;
				18'b010110010000100010: oled_data = 16'b1001000101100111;
				18'b010110010010100010: oled_data = 16'b1000100101000110;
				18'b010110010100100010: oled_data = 16'b1010101000001000;
				18'b010110010110100010: oled_data = 16'b1011001001001001;
				18'b010110011000100010: oled_data = 16'b1011001001001001;
				18'b010110011010100010: oled_data = 16'b1011001001001001;
				18'b010110011100100010: oled_data = 16'b1011001001001001;
				18'b010110011110100010: oled_data = 16'b1011001001001001;
				18'b010110100000100010: oled_data = 16'b1011001000101001;
				18'b010110100010100010: oled_data = 16'b1011001000101000;
				18'b010110100100100010: oled_data = 16'b1011001000001000;
				18'b010110100110100010: oled_data = 16'b1010101000001000;
				18'b010100011000100011: oled_data = 16'b1101110011110110;
				18'b010100011010100011: oled_data = 16'b1101110011010110;
				18'b010100011100100011: oled_data = 16'b1101110011110110;
				18'b010100011110100011: oled_data = 16'b1101110011010110;
				18'b010100100000100011: oled_data = 16'b1110010011010110;
				18'b010100100010100011: oled_data = 16'b1101110010010101;
				18'b010100100100100011: oled_data = 16'b1100110000110011;
				18'b010100100110100011: oled_data = 16'b1101110010110101;
				18'b010100101000100011: oled_data = 16'b1101010001110100;
				18'b010100101010100011: oled_data = 16'b1101110011010101;
				18'b010100101100100011: oled_data = 16'b1101010001110100;
				18'b010100101110100011: oled_data = 16'b1101110011010101;
				18'b010100110000100011: oled_data = 16'b1101110011010101;
				18'b010100110010100011: oled_data = 16'b1101110011010101;
				18'b010100110100100011: oled_data = 16'b1101110011010101;
				18'b010100110110100011: oled_data = 16'b1101110011010101;
				18'b010100111000100011: oled_data = 16'b1110010011010101;
				18'b010100111010100011: oled_data = 16'b1101010001010100;
				18'b010100111100100011: oled_data = 16'b1101010100110110;
				18'b010100111110100011: oled_data = 16'b1110011001111010;
				18'b010101000000100011: oled_data = 16'b1101110010110101;
				18'b010101000010100011: oled_data = 16'b1101110101110111;
				18'b010101000100100011: oled_data = 16'b1110111100011011;
				18'b010101000110100011: oled_data = 16'b1110111100011010;
				18'b010101001000100011: oled_data = 16'b1110111100111011;
				18'b010101001010100011: oled_data = 16'b1110111101011011;
				18'b010101001100100011: oled_data = 16'b1110111101011011;
				18'b010101001110100011: oled_data = 16'b1101011000110111;
				18'b010101010000100011: oled_data = 16'b1110011011011010;
				18'b010101010010100011: oled_data = 16'b1110111100011011;
				18'b010101010100100011: oled_data = 16'b1110111010011010;
				18'b010101010110100011: oled_data = 16'b1101110011110110;
				18'b010101011000100011: oled_data = 16'b1110010011010110;
				18'b010101011010100011: oled_data = 16'b1110010011010110;
				18'b010101011100100011: oled_data = 16'b1110010011010110;
				18'b010101011110100011: oled_data = 16'b1101110010110101;
				18'b010101100000100011: oled_data = 16'b1101010001110100;
				18'b010101100010100011: oled_data = 16'b1101010101010110;
				18'b010101100100100011: oled_data = 16'b1110011100011010;
				18'b010101100110100011: oled_data = 16'b1110011100011010;
				18'b010101101000100011: oled_data = 16'b1110111100011010;
				18'b010101101010100011: oled_data = 16'b1110011100011010;
				18'b010101101100100011: oled_data = 16'b1110011100011010;
				18'b010101101110100011: oled_data = 16'b1110111100011010;
				18'b010101110000100011: oled_data = 16'b1110111100011010;
				18'b010101110010100011: oled_data = 16'b1110111100011010;
				18'b010101110100100011: oled_data = 16'b1110111100011010;
				18'b010101110110100011: oled_data = 16'b1110011011111010;
				18'b010101111000100011: oled_data = 16'b1101111010111001;
				18'b010101111010100011: oled_data = 16'b1110111100111011;
				18'b010101111100100011: oled_data = 16'b1101110110010110;
				18'b010101111110100011: oled_data = 16'b1110010100010100;
				18'b010110000000100011: oled_data = 16'b1100001100101100;
				18'b010110000010100011: oled_data = 16'b1011001000101000;
				18'b010110000100100011: oled_data = 16'b1011101001001001;
				18'b010110000110100011: oled_data = 16'b1011001001001001;
				18'b010110001000100011: oled_data = 16'b1011001001001001;
				18'b010110001010100011: oled_data = 16'b1011001000101001;
				18'b010110001100100011: oled_data = 16'b1010101000101001;
				18'b010110001110100011: oled_data = 16'b1010000111101000;
				18'b010110010000100011: oled_data = 16'b1000100101000110;
				18'b010110010010100011: oled_data = 16'b1001100111001000;
				18'b010110010100100011: oled_data = 16'b1011001001001001;
				18'b010110010110100011: oled_data = 16'b1011001001001001;
				18'b010110011000100011: oled_data = 16'b1011001001001001;
				18'b010110011010100011: oled_data = 16'b1011001001001001;
				18'b010110011100100011: oled_data = 16'b1011001000101001;
				18'b010110011110100011: oled_data = 16'b1011001000101001;
				18'b010110100000100011: oled_data = 16'b1011001000101001;
				18'b010110100010100011: oled_data = 16'b1011001000101000;
				18'b010110100100100011: oled_data = 16'b1011001000001000;
				18'b010110100110100011: oled_data = 16'b1010101000001000;
				18'b010100011000100100: oled_data = 16'b1101110011010110;
				18'b010100011010100100: oled_data = 16'b1101110011010110;
				18'b010100011100100100: oled_data = 16'b1101110011110110;
				18'b010100011110100100: oled_data = 16'b1101110011110110;
				18'b010100100000100100: oled_data = 16'b1110010011110110;
				18'b010100100010100100: oled_data = 16'b1101010001010011;
				18'b010100100100100100: oled_data = 16'b1101010001010100;
				18'b010100100110100100: oled_data = 16'b1101110010010101;
				18'b010100101000100100: oled_data = 16'b1101010010010101;
				18'b010100101010100100: oled_data = 16'b1101110010110101;
				18'b010100101100100100: oled_data = 16'b1101010010010100;
				18'b010100101110100100: oled_data = 16'b1101110011010110;
				18'b010100110000100100: oled_data = 16'b1101110011010101;
				18'b010100110010100100: oled_data = 16'b1101110011010101;
				18'b010100110100100100: oled_data = 16'b1101110011010101;
				18'b010100110110100100: oled_data = 16'b1101110011010101;
				18'b010100111000100100: oled_data = 16'b1101110011010110;
				18'b010100111010100100: oled_data = 16'b1101010001010100;
				18'b010100111100100100: oled_data = 16'b1101110110010111;
				18'b010100111110100100: oled_data = 16'b1110111001111010;
				18'b010101000000100100: oled_data = 16'b1101110011110101;
				18'b010101000010100100: oled_data = 16'b1110111010011001;
				18'b010101000100100100: oled_data = 16'b1110111100011010;
				18'b010101000110100100: oled_data = 16'b1110011011111010;
				18'b010101001000100100: oled_data = 16'b1011010101110100;
				18'b010101001010100100: oled_data = 16'b1010010100010011;
				18'b010101001100100100: oled_data = 16'b1011010110010101;
				18'b010101001110100100: oled_data = 16'b1011110110110101;
				18'b010101010000100100: oled_data = 16'b1100010111110111;
				18'b010101010010100100: oled_data = 16'b1101011000111000;
				18'b010101010100100100: oled_data = 16'b1100110111110111;
				18'b010101010110100100: oled_data = 16'b1100010010010011;
				18'b010101011000100100: oled_data = 16'b1101010010010100;
				18'b010101011010100100: oled_data = 16'b1101010010110100;
				18'b010101011100100100: oled_data = 16'b1101010010110101;
				18'b010101011110100100: oled_data = 16'b1101010010010100;
				18'b010101100000100100: oled_data = 16'b1100110011010101;
				18'b010101100010100100: oled_data = 16'b1110011010011010;
				18'b010101100100100100: oled_data = 16'b1110111100111011;
				18'b010101100110100100: oled_data = 16'b1110011100011011;
				18'b010101101000100100: oled_data = 16'b1110111100011010;
				18'b010101101010100100: oled_data = 16'b1110111100011010;
				18'b010101101100100100: oled_data = 16'b1110111100011010;
				18'b010101101110100100: oled_data = 16'b1110111100011010;
				18'b010101110000100100: oled_data = 16'b1110011100011010;
				18'b010101110010100100: oled_data = 16'b1110111100011010;
				18'b010101110100100100: oled_data = 16'b1110111100011011;
				18'b010101110110100100: oled_data = 16'b1101111010111010;
				18'b010101111000100100: oled_data = 16'b1110111100011010;
				18'b010101111010100100: oled_data = 16'b1110011011111010;
				18'b010101111100100100: oled_data = 16'b1101110100110101;
				18'b010101111110100100: oled_data = 16'b1110110011110011;
				18'b010110000000100100: oled_data = 16'b1011001010101011;
				18'b010110000010100100: oled_data = 16'b1011001000101001;
				18'b010110000100100100: oled_data = 16'b1011001001001001;
				18'b010110000110100100: oled_data = 16'b1011001001001001;
				18'b010110001000100100: oled_data = 16'b1011001001001001;
				18'b010110001010100100: oled_data = 16'b1010101000101000;
				18'b010110001100100100: oled_data = 16'b1011001000101001;
				18'b010110001110100100: oled_data = 16'b1001000101100110;
				18'b010110010000100100: oled_data = 16'b1001000101100111;
				18'b010110010010100100: oled_data = 16'b1011001000101001;
				18'b010110010100100100: oled_data = 16'b1011001001001001;
				18'b010110010110100100: oled_data = 16'b1011001000101001;
				18'b010110011000100100: oled_data = 16'b1011001001001001;
				18'b010110011010100100: oled_data = 16'b1011001001001001;
				18'b010110011100100100: oled_data = 16'b1011001001001001;
				18'b010110011110100100: oled_data = 16'b1011001001001001;
				18'b010110100000100100: oled_data = 16'b1011001000101001;
				18'b010110100010100100: oled_data = 16'b1011001000101000;
				18'b010110100100100100: oled_data = 16'b1010101000101000;
				18'b010110100110100100: oled_data = 16'b1010101000101000;
				18'b010100011000100101: oled_data = 16'b1101110011010110;
				18'b010100011010100101: oled_data = 16'b1101110011010110;
				18'b010100011100100101: oled_data = 16'b1101110011010110;
				18'b010100011110100101: oled_data = 16'b1101110011010110;
				18'b010100100000100101: oled_data = 16'b1110010011110110;
				18'b010100100010100101: oled_data = 16'b1101010001010100;
				18'b010100100100100101: oled_data = 16'b1101110010110101;
				18'b010100100110100101: oled_data = 16'b1100110000110011;
				18'b010100101000100101: oled_data = 16'b1101110010110101;
				18'b010100101010100101: oled_data = 16'b1101010010010100;
				18'b010100101100100101: oled_data = 16'b1101010010010101;
				18'b010100101110100101: oled_data = 16'b1101110011010110;
				18'b010100110000100101: oled_data = 16'b1101110011010101;
				18'b010100110010100101: oled_data = 16'b1101110011010101;
				18'b010100110100100101: oled_data = 16'b1101110011010101;
				18'b010100110110100101: oled_data = 16'b1101110011010101;
				18'b010100111000100101: oled_data = 16'b1101110011010101;
				18'b010100111010100101: oled_data = 16'b1101010001110100;
				18'b010100111100100101: oled_data = 16'b1101110111111000;
				18'b010100111110100101: oled_data = 16'b1110011001111001;
				18'b010101000000100101: oled_data = 16'b1101110111010111;
				18'b010101000010100101: oled_data = 16'b1110111100011010;
				18'b010101000100100101: oled_data = 16'b1110111100011010;
				18'b010101000110100101: oled_data = 16'b1100111000110111;
				18'b010101001000100101: oled_data = 16'b0101001001101000;
				18'b010101001010100101: oled_data = 16'b0010100100100100;
				18'b010101001100100101: oled_data = 16'b0011000101000100;
				18'b010101001110100101: oled_data = 16'b0011000101100100;
				18'b010101010000100101: oled_data = 16'b0011000110000101;
				18'b010101010010100101: oled_data = 16'b0011100110000110;
				18'b010101010100100101: oled_data = 16'b0011100110000110;
				18'b010101010110100101: oled_data = 16'b0101100111001000;
				18'b010101011000100101: oled_data = 16'b0110101000101010;
				18'b010101011010100101: oled_data = 16'b0111001000101010;
				18'b010101011100100101: oled_data = 16'b0111001000101010;
				18'b010101011110100101: oled_data = 16'b1100010001110011;
				18'b010101100000100101: oled_data = 16'b1101111001011001;
				18'b010101100010100101: oled_data = 16'b1110111100011011;
				18'b010101100100100101: oled_data = 16'b1110111100011011;
				18'b010101100110100101: oled_data = 16'b1110111100011011;
				18'b010101101000100101: oled_data = 16'b1110111100011010;
				18'b010101101010100101: oled_data = 16'b1110111100011010;
				18'b010101101100100101: oled_data = 16'b1110111100011010;
				18'b010101101110100101: oled_data = 16'b1110111100011010;
				18'b010101110000100101: oled_data = 16'b1110111100011010;
				18'b010101110010100101: oled_data = 16'b1110111100011010;
				18'b010101110100100101: oled_data = 16'b1101111010111001;
				18'b010101110110100101: oled_data = 16'b1110011011011010;
				18'b010101111000100101: oled_data = 16'b1110111100111011;
				18'b010101111010100101: oled_data = 16'b1110011010011010;
				18'b010101111100100101: oled_data = 16'b1101110011110100;
				18'b010101111110100101: oled_data = 16'b1110010011010011;
				18'b010110000000100101: oled_data = 16'b1011001001101001;
				18'b010110000010100101: oled_data = 16'b1011001001001001;
				18'b010110000100100101: oled_data = 16'b1011001001001001;
				18'b010110000110100101: oled_data = 16'b1011001001001001;
				18'b010110001000100101: oled_data = 16'b1011101010101010;
				18'b010110001010100101: oled_data = 16'b1011001010001001;
				18'b010110001100100101: oled_data = 16'b1010000111100111;
				18'b010110001110100101: oled_data = 16'b1000100101000110;
				18'b010110010000100101: oled_data = 16'b1010000111101001;
				18'b010110010010100101: oled_data = 16'b1011001001001001;
				18'b010110010100100101: oled_data = 16'b1011001000101000;
				18'b010110010110100101: oled_data = 16'b1011101110101111;
				18'b010110011000100101: oled_data = 16'b1011001010101011;
				18'b010110011010100101: oled_data = 16'b1011001001001001;
				18'b010110011100100101: oled_data = 16'b1011101010001010;
				18'b010110011110100101: oled_data = 16'b1011001001001001;
				18'b010110100000100101: oled_data = 16'b1011001000101001;
				18'b010110100010100101: oled_data = 16'b1011001000101000;
				18'b010110100100100101: oled_data = 16'b1010101000101000;
				18'b010110100110100101: oled_data = 16'b1010101000101000;
				18'b010100011000100110: oled_data = 16'b1101110011010110;
				18'b010100011010100110: oled_data = 16'b1101110011010110;
				18'b010100011100100110: oled_data = 16'b1110010010110101;
				18'b010100011110100110: oled_data = 16'b1110010010110101;
				18'b010100100000100110: oled_data = 16'b1101110011010101;
				18'b010100100010100110: oled_data = 16'b1101010001110100;
				18'b010100100100100110: oled_data = 16'b1101110010010101;
				18'b010100100110100110: oled_data = 16'b1100001111110010;
				18'b010100101000100110: oled_data = 16'b1101110011010110;
				18'b010100101010100110: oled_data = 16'b1100110000110011;
				18'b010100101100100110: oled_data = 16'b1101110010110101;
				18'b010100101110100110: oled_data = 16'b1101110011010110;
				18'b010100110000100110: oled_data = 16'b1101110011010101;
				18'b010100110010100110: oled_data = 16'b1101110011010101;
				18'b010100110100100110: oled_data = 16'b1101110011010101;
				18'b010100110110100110: oled_data = 16'b1101110011010101;
				18'b010100111000100110: oled_data = 16'b1101110010110101;
				18'b010100111010100110: oled_data = 16'b1101010001110100;
				18'b010100111100100110: oled_data = 16'b1110011001011001;
				18'b010100111110100110: oled_data = 16'b1110011011111010;
				18'b010101000000100110: oled_data = 16'b1110011011111010;
				18'b010101000010100110: oled_data = 16'b1110111100011010;
				18'b010101000100100110: oled_data = 16'b1110111100011010;
				18'b010101000110100110: oled_data = 16'b1101011001111000;
				18'b010101001000100110: oled_data = 16'b1010010011110011;
				18'b010101001010100110: oled_data = 16'b1000001111101111;
				18'b010101001100100110: oled_data = 16'b0110101100101100;
				18'b010101001110100110: oled_data = 16'b0101101010101010;
				18'b010101010000100110: oled_data = 16'b0101101010001001;
				18'b010101010010100110: oled_data = 16'b0101001001001000;
				18'b010101010100100110: oled_data = 16'b0101001000101000;
				18'b010101010110100110: oled_data = 16'b0110001001001001;
				18'b010101011000100110: oled_data = 16'b0101101000001000;
				18'b010101011010100110: oled_data = 16'b0100100110000110;
				18'b010101011100100110: oled_data = 16'b0111001010101011;
				18'b010101011110100110: oled_data = 16'b1101111000011000;
				18'b010101100000100110: oled_data = 16'b1110111100011011;
				18'b010101100010100110: oled_data = 16'b1110111100011010;
				18'b010101100100100110: oled_data = 16'b1110111100011010;
				18'b010101100110100110: oled_data = 16'b1110111100011010;
				18'b010101101000100110: oled_data = 16'b1110111100011010;
				18'b010101101010100110: oled_data = 16'b1110111100011010;
				18'b010101101100100110: oled_data = 16'b1110111100011010;
				18'b010101101110100110: oled_data = 16'b1110111100011010;
				18'b010101110000100110: oled_data = 16'b1110111100011010;
				18'b010101110010100110: oled_data = 16'b1110011011111010;
				18'b010101110100100110: oled_data = 16'b1101111010011001;
				18'b010101110110100110: oled_data = 16'b1110111100011011;
				18'b010101111000100110: oled_data = 16'b1110111100111011;
				18'b010101111010100110: oled_data = 16'b1100010100110101;
				18'b010101111100100110: oled_data = 16'b1100110001110010;
				18'b010101111110100110: oled_data = 16'b1101110001110001;
				18'b010110000000100110: oled_data = 16'b1010101000101001;
				18'b010110000010100110: oled_data = 16'b1011001001001001;
				18'b010110000100100110: oled_data = 16'b1011001010101010;
				18'b010110000110100110: oled_data = 16'b1101010000110000;
				18'b010110001000100110: oled_data = 16'b1110010010110011;
				18'b010110001010100110: oled_data = 16'b1100101110101111;
				18'b010110001100100110: oled_data = 16'b1010000111101000;
				18'b010110001110100110: oled_data = 16'b1001100110000111;
				18'b010110010000100110: oled_data = 16'b1011001001101010;
				18'b010110010010100110: oled_data = 16'b1011001001001001;
				18'b010110010100100110: oled_data = 16'b1011001001101010;
				18'b010110010110100110: oled_data = 16'b1100011000111001;
				18'b010110011000100110: oled_data = 16'b1011001111110000;
				18'b010110011010100110: oled_data = 16'b1011001000001000;
				18'b010110011100100110: oled_data = 16'b1011001001001001;
				18'b010110011110100110: oled_data = 16'b1011001000101001;
				18'b010110100000100110: oled_data = 16'b1011001000101001;
				18'b010110100010100110: oled_data = 16'b1011001000101000;
				18'b010110100100100110: oled_data = 16'b1010101000101000;
				18'b010110100110100110: oled_data = 16'b1010101000101000;
				18'b010100011000100111: oled_data = 16'b1101110011010110;
				18'b010100011010100111: oled_data = 16'b1101110011010110;
				18'b010100011100100111: oled_data = 16'b1110010010110101;
				18'b010100011110100111: oled_data = 16'b1110010011010101;
				18'b010100100000100111: oled_data = 16'b1101110010110101;
				18'b010100100010100111: oled_data = 16'b1101010010010101;
				18'b010100100100100111: oled_data = 16'b1100110000110011;
				18'b010100100110100111: oled_data = 16'b1100001111110010;
				18'b010100101000100111: oled_data = 16'b1101110011010110;
				18'b010100101010100111: oled_data = 16'b1100001111110010;
				18'b010100101100100111: oled_data = 16'b1101110011010101;
				18'b010100101110100111: oled_data = 16'b1110010011010110;
				18'b010100110000100111: oled_data = 16'b1110010011010110;
				18'b010100110010100111: oled_data = 16'b1110010011010110;
				18'b010100110100100111: oled_data = 16'b1110010011010110;
				18'b010100110110100111: oled_data = 16'b1110010011110110;
				18'b010100111000100111: oled_data = 16'b1101110010110101;
				18'b010100111010100111: oled_data = 16'b1101010010010100;
				18'b010100111100100111: oled_data = 16'b1110011010111010;
				18'b010100111110100111: oled_data = 16'b1110111100011010;
				18'b010101000000100111: oled_data = 16'b1110111100011010;
				18'b010101000010100111: oled_data = 16'b1110111100011010;
				18'b010101000100100111: oled_data = 16'b1110111100011010;
				18'b010101000110100111: oled_data = 16'b1110111100011011;
				18'b010101001000100111: oled_data = 16'b1110111100111100;
				18'b010101001010100111: oled_data = 16'b1110111100111011;
				18'b010101001100100111: oled_data = 16'b1110111100011010;
				18'b010101001110100111: oled_data = 16'b1110011100011010;
				18'b010101010000100111: oled_data = 16'b1110011011111010;
				18'b010101010010100111: oled_data = 16'b1101111011011010;
				18'b010101010100100111: oled_data = 16'b1110011011011010;
				18'b010101010110100111: oled_data = 16'b1011010011010010;
				18'b010101011000100111: oled_data = 16'b0101101000001000;
				18'b010101011010100111: oled_data = 16'b0101000111100111;
				18'b010101011100100111: oled_data = 16'b1100010110010110;
				18'b010101011110100111: oled_data = 16'b1110111011111011;
				18'b010101100000100111: oled_data = 16'b1110011100011010;
				18'b010101100010100111: oled_data = 16'b1110111100011010;
				18'b010101100100100111: oled_data = 16'b1110111100011010;
				18'b010101100110100111: oled_data = 16'b1110111100011010;
				18'b010101101000100111: oled_data = 16'b1110111100011010;
				18'b010101101010100111: oled_data = 16'b1110111100011010;
				18'b010101101100100111: oled_data = 16'b1110111100011010;
				18'b010101101110100111: oled_data = 16'b1110111100011010;
				18'b010101110000100111: oled_data = 16'b1110011100011010;
				18'b010101110010100111: oled_data = 16'b1101111010011000;
				18'b010101110100100111: oled_data = 16'b1110011011111010;
				18'b010101110110100111: oled_data = 16'b1110111100111011;
				18'b010101111000100111: oled_data = 16'b1101111000111000;
				18'b010101111010100111: oled_data = 16'b1010101111110001;
				18'b010101111100100111: oled_data = 16'b1101010010110011;
				18'b010101111110100111: oled_data = 16'b1101010000110000;
				18'b010110000000100111: oled_data = 16'b1010101000101000;
				18'b010110000010100111: oled_data = 16'b1011001001001001;
				18'b010110000100100111: oled_data = 16'b1101010001010001;
				18'b010110000110100111: oled_data = 16'b1110110011110011;
				18'b010110001000100111: oled_data = 16'b1100001100001101;
				18'b010110001010100111: oled_data = 16'b1011001000101001;
				18'b010110001100100111: oled_data = 16'b1011001000101001;
				18'b010110001110100111: oled_data = 16'b1011001001001001;
				18'b010110010000100111: oled_data = 16'b1011001001101010;
				18'b010110010010100111: oled_data = 16'b1011001000101001;
				18'b010110010100100111: oled_data = 16'b1011101111110000;
				18'b010110010110100111: oled_data = 16'b1011111100011100;
				18'b010110011000100111: oled_data = 16'b1011110111010111;
				18'b010110011010100111: oled_data = 16'b1011001001001001;
				18'b010110011100100111: oled_data = 16'b1011001000101001;
				18'b010110011110100111: oled_data = 16'b1011001001001001;
				18'b010110100000100111: oled_data = 16'b1011001000101000;
				18'b010110100010100111: oled_data = 16'b1010101000001000;
				18'b010110100100100111: oled_data = 16'b1010000111101000;
				18'b010110100110100111: oled_data = 16'b1010101000001000;
				18'b010100011000101000: oled_data = 16'b1101110011010101;
				18'b010100011010101000: oled_data = 16'b1101110011010101;
				18'b010100011100101000: oled_data = 16'b1101110011010101;
				18'b010100011110101000: oled_data = 16'b1101110011010110;
				18'b010100100000101000: oled_data = 16'b1101010001110100;
				18'b010100100010101000: oled_data = 16'b1101010010010100;
				18'b010100100100101000: oled_data = 16'b1011101110110001;
				18'b010100100110101000: oled_data = 16'b1100110000010011;
				18'b010100101000101000: oled_data = 16'b1101110010110101;
				18'b010100101010101000: oled_data = 16'b1100001111110010;
				18'b010100101100101000: oled_data = 16'b1101110011010110;
				18'b010100101110101000: oled_data = 16'b1101110011010101;
				18'b010100110000101000: oled_data = 16'b1101110011010101;
				18'b010100110010101000: oled_data = 16'b1101110011010101;
				18'b010100110100101000: oled_data = 16'b1101110011010110;
				18'b010100110110101000: oled_data = 16'b1110010011110110;
				18'b010100111000101000: oled_data = 16'b1101010010110101;
				18'b010100111010101000: oled_data = 16'b1100110010110100;
				18'b010100111100101000: oled_data = 16'b1110011011011010;
				18'b010100111110101000: oled_data = 16'b1110011100011010;
				18'b010101000000101000: oled_data = 16'b1110111100011010;
				18'b010101000010101000: oled_data = 16'b1110111100011010;
				18'b010101000100101000: oled_data = 16'b1110111100011010;
				18'b010101000110101000: oled_data = 16'b1110111100011010;
				18'b010101001000101000: oled_data = 16'b1110111100011011;
				18'b010101001010101000: oled_data = 16'b1110111100011010;
				18'b010101001100101000: oled_data = 16'b1110111100011010;
				18'b010101001110101000: oled_data = 16'b1110111100011010;
				18'b010101010000101000: oled_data = 16'b1110011100011010;
				18'b010101010010101000: oled_data = 16'b1110111100111011;
				18'b010101010100101000: oled_data = 16'b1110011010011001;
				18'b010101010110101000: oled_data = 16'b0111001010101011;
				18'b010101011000101000: oled_data = 16'b0100100110100111;
				18'b010101011010101000: oled_data = 16'b1011010100110100;
				18'b010101011100101000: oled_data = 16'b1111011100111011;
				18'b010101011110101000: oled_data = 16'b1110111100011010;
				18'b010101100000101000: oled_data = 16'b1110111100011010;
				18'b010101100010101000: oled_data = 16'b1110111100011010;
				18'b010101100100101000: oled_data = 16'b1110111100011010;
				18'b010101100110101000: oled_data = 16'b1110111100011010;
				18'b010101101000101000: oled_data = 16'b1110111100011010;
				18'b010101101010101000: oled_data = 16'b1110111100011010;
				18'b010101101100101000: oled_data = 16'b1110111100011010;
				18'b010101101110101000: oled_data = 16'b1110111100011010;
				18'b010101110000101000: oled_data = 16'b1101111010111001;
				18'b010101110010101000: oled_data = 16'b1110011011111010;
				18'b010101110100101000: oled_data = 16'b1110111100011011;
				18'b010101110110101000: oled_data = 16'b1101111001111000;
				18'b010101111000101000: oled_data = 16'b1100110101010101;
				18'b010101111010101000: oled_data = 16'b1101110101110110;
				18'b010101111100101000: oled_data = 16'b1101110100010100;
				18'b010101111110101000: oled_data = 16'b1100101111001111;
				18'b010110000000101000: oled_data = 16'b1010101000001000;
				18'b010110000010101000: oled_data = 16'b1011101011101100;
				18'b010110000100101000: oled_data = 16'b1110110011110100;
				18'b010110000110101000: oled_data = 16'b1100101101101110;
				18'b010110001000101000: oled_data = 16'b1011001000101001;
				18'b010110001010101000: oled_data = 16'b1011001001001001;
				18'b010110001100101000: oled_data = 16'b1011001001001001;
				18'b010110001110101000: oled_data = 16'b1011001001001001;
				18'b010110010000101000: oled_data = 16'b1011001001001001;
				18'b010110010010101000: oled_data = 16'b1011001001001001;
				18'b010110010100101000: oled_data = 16'b1100010110110110;
				18'b010110010110101000: oled_data = 16'b1011111100011100;
				18'b010110011000101000: oled_data = 16'b1011111011111011;
				18'b010110011010101000: oled_data = 16'b1011001101101110;
				18'b010110011100101000: oled_data = 16'b1010101000001000;
				18'b010110011110101000: oled_data = 16'b1010101000001000;
				18'b010110100000101000: oled_data = 16'b1010001000001000;
				18'b010110100010101000: oled_data = 16'b1010001000001000;
				18'b010110100100101000: oled_data = 16'b1010101000001000;
				18'b010110100110101000: oled_data = 16'b1010101000001000;
				18'b010100011000101001: oled_data = 16'b1101110011010101;
				18'b010100011010101001: oled_data = 16'b1101110011010101;
				18'b010100011100101001: oled_data = 16'b1101110011010101;
				18'b010100011110101001: oled_data = 16'b1101110011010101;
				18'b010100100000101001: oled_data = 16'b1101110010010101;
				18'b010100100010101001: oled_data = 16'b1100110001010100;
				18'b010100100100101001: oled_data = 16'b1011001101110001;
				18'b010100100110101001: oled_data = 16'b1100110001010011;
				18'b010100101000101001: oled_data = 16'b1101010010010100;
				18'b010100101010101001: oled_data = 16'b1100001111110010;
				18'b010100101100101001: oled_data = 16'b1110010011010110;
				18'b010100101110101001: oled_data = 16'b1101110011010101;
				18'b010100110000101001: oled_data = 16'b1101110011010110;
				18'b010100110010101001: oled_data = 16'b1110010011010110;
				18'b010100110100101001: oled_data = 16'b1110010011010110;
				18'b010100110110101001: oled_data = 16'b1110010011110110;
				18'b010100111000101001: oled_data = 16'b1101110010010101;
				18'b010100111010101001: oled_data = 16'b1101010011010101;
				18'b010100111100101001: oled_data = 16'b1110111011111010;
				18'b010100111110101001: oled_data = 16'b1110011100011010;
				18'b010101000000101001: oled_data = 16'b1110111100011010;
				18'b010101000010101001: oled_data = 16'b1110111100011010;
				18'b010101000100101001: oled_data = 16'b1110111100011010;
				18'b010101000110101001: oled_data = 16'b1110111100011010;
				18'b010101001000101001: oled_data = 16'b1110111100011010;
				18'b010101001010101001: oled_data = 16'b1110111100011010;
				18'b010101001100101001: oled_data = 16'b1110111100011010;
				18'b010101001110101001: oled_data = 16'b1110111100011010;
				18'b010101010000101001: oled_data = 16'b1110111100011011;
				18'b010101010010101001: oled_data = 16'b1110011011111010;
				18'b010101010100101001: oled_data = 16'b0111101101001101;
				18'b010101010110101001: oled_data = 16'b0011100100100101;
				18'b010101011000101001: oled_data = 16'b1001010000110000;
				18'b010101011010101001: oled_data = 16'b1110111100111011;
				18'b010101011100101001: oled_data = 16'b1110111100011010;
				18'b010101011110101001: oled_data = 16'b1110111100011010;
				18'b010101100000101001: oled_data = 16'b1110111100011010;
				18'b010101100010101001: oled_data = 16'b1110111100011010;
				18'b010101100100101001: oled_data = 16'b1110111100011010;
				18'b010101100110101001: oled_data = 16'b1110111100011010;
				18'b010101101000101001: oled_data = 16'b1110111100011010;
				18'b010101101010101001: oled_data = 16'b1110111100011010;
				18'b010101101100101001: oled_data = 16'b1110111100011010;
				18'b010101101110101001: oled_data = 16'b1101111010111001;
				18'b010101110000101001: oled_data = 16'b1101111011011001;
				18'b010101110010101001: oled_data = 16'b1110111100111011;
				18'b010101110100101001: oled_data = 16'b1101111010011001;
				18'b010101110110101001: oled_data = 16'b1101010111010110;
				18'b010101111000101001: oled_data = 16'b1110111010111001;
				18'b010101111010101001: oled_data = 16'b1110011011011010;
				18'b010101111100101001: oled_data = 16'b1101110100110100;
				18'b010101111110101001: oled_data = 16'b1100101110001110;
				18'b010110000000101001: oled_data = 16'b1011001000001000;
				18'b010110000010101001: oled_data = 16'b1100101110101110;
				18'b010110000100101001: oled_data = 16'b1110010011010010;
				18'b010110000110101001: oled_data = 16'b1011101010001010;
				18'b010110001000101001: oled_data = 16'b1011001001001001;
				18'b010110001010101001: oled_data = 16'b1011001001001001;
				18'b010110001100101001: oled_data = 16'b1011001001001001;
				18'b010110001110101001: oled_data = 16'b1011001001001001;
				18'b010110010000101001: oled_data = 16'b1011001000101001;
				18'b010110010010101001: oled_data = 16'b1011001101101110;
				18'b010110010100101001: oled_data = 16'b1100011011011011;
				18'b010110010110101001: oled_data = 16'b1011111011111011;
				18'b010110011000101001: oled_data = 16'b1011111100011100;
				18'b010110011010101001: oled_data = 16'b1011110101010101;
				18'b010110011100101001: oled_data = 16'b1010101000101001;
				18'b010110011110101001: oled_data = 16'b1011001000101000;
				18'b010110100000101001: oled_data = 16'b1011001000101000;
				18'b010110100010101001: oled_data = 16'b1010101000101000;
				18'b010110100100101001: oled_data = 16'b1010101000001000;
				18'b010110100110101001: oled_data = 16'b1010101000001000;
				18'b010100011000101010: oled_data = 16'b1101110011010101;
				18'b010100011010101010: oled_data = 16'b1101110011010101;
				18'b010100011100101010: oled_data = 16'b1101110011010101;
				18'b010100011110101010: oled_data = 16'b1101110010110101;
				18'b010100100000101010: oled_data = 16'b1101010010010100;
				18'b010100100010101010: oled_data = 16'b1100001111110010;
				18'b010100100100101010: oled_data = 16'b1011001101110000;
				18'b010100100110101010: oled_data = 16'b1101010001110100;
				18'b010100101000101010: oled_data = 16'b1101010010010100;
				18'b010100101010101010: oled_data = 16'b1100010000010010;
				18'b010100101100101010: oled_data = 16'b1110010011010110;
				18'b010100101110101010: oled_data = 16'b1110010011010110;
				18'b010100110000101010: oled_data = 16'b1110010011010110;
				18'b010100110010101010: oled_data = 16'b1110010011010110;
				18'b010100110100101010: oled_data = 16'b1110010011010110;
				18'b010100110110101010: oled_data = 16'b1110010011110110;
				18'b010100111000101010: oled_data = 16'b1101110010010101;
				18'b010100111010101010: oled_data = 16'b1101010100010101;
				18'b010100111100101010: oled_data = 16'b1110011011111010;
				18'b010100111110101010: oled_data = 16'b1110111100011010;
				18'b010101000000101010: oled_data = 16'b1110111100011010;
				18'b010101000010101010: oled_data = 16'b1110111100011010;
				18'b010101000100101010: oled_data = 16'b1110111100011010;
				18'b010101000110101010: oled_data = 16'b1110111100011010;
				18'b010101001000101010: oled_data = 16'b1110111100011010;
				18'b010101001010101010: oled_data = 16'b1110111100011010;
				18'b010101001100101010: oled_data = 16'b1110111100011010;
				18'b010101001110101010: oled_data = 16'b1110111100011011;
				18'b010101010000101010: oled_data = 16'b1110111100111011;
				18'b010101010010101010: oled_data = 16'b1000001111001110;
				18'b010101010100101010: oled_data = 16'b0011000100100100;
				18'b010101010110101010: oled_data = 16'b0111001101001101;
				18'b010101011000101010: oled_data = 16'b1110011011111011;
				18'b010101011010101010: oled_data = 16'b1110111100011011;
				18'b010101011100101010: oled_data = 16'b1110111100011010;
				18'b010101011110101010: oled_data = 16'b1110111100011010;
				18'b010101100000101010: oled_data = 16'b1110111100011010;
				18'b010101100010101010: oled_data = 16'b1110111100011010;
				18'b010101100100101010: oled_data = 16'b1110111100011010;
				18'b010101100110101010: oled_data = 16'b1110111100011010;
				18'b010101101000101010: oled_data = 16'b1110111100011010;
				18'b010101101010101010: oled_data = 16'b1110111100011010;
				18'b010101101100101010: oled_data = 16'b1110111100011010;
				18'b010101101110101010: oled_data = 16'b1110011011111010;
				18'b010101110000101010: oled_data = 16'b1110111100111010;
				18'b010101110010101010: oled_data = 16'b1101111010111001;
				18'b010101110100101010: oled_data = 16'b1101111001011000;
				18'b010101110110101010: oled_data = 16'b1110111011111010;
				18'b010101111000101010: oled_data = 16'b1110111100011011;
				18'b010101111010101010: oled_data = 16'b1110011011011010;
				18'b010101111100101010: oled_data = 16'b1101010100110100;
				18'b010101111110101010: oled_data = 16'b1100001101001101;
				18'b010110000000101010: oled_data = 16'b1010101000001000;
				18'b010110000010101010: oled_data = 16'b1101010000110000;
				18'b010110000100101010: oled_data = 16'b1101110000010000;
				18'b010110000110101010: oled_data = 16'b1011001001001001;
				18'b010110001000101010: oled_data = 16'b1011101001001001;
				18'b010110001010101010: oled_data = 16'b1011001001001001;
				18'b010110001100101010: oled_data = 16'b1011001001001001;
				18'b010110001110101010: oled_data = 16'b1011001001001001;
				18'b010110010000101010: oled_data = 16'b1011001000101001;
				18'b010110010010101010: oled_data = 16'b1011110101110110;
				18'b010110010100101010: oled_data = 16'b1011111100011100;
				18'b010110010110101010: oled_data = 16'b1011111011111011;
				18'b010110011000101010: oled_data = 16'b1011111011111100;
				18'b010110011010101010: oled_data = 16'b1100011010111011;
				18'b010110011100101010: oled_data = 16'b1011001100001100;
				18'b010110011110101010: oled_data = 16'b1010101000101000;
				18'b010110100000101010: oled_data = 16'b1011001000101001;
				18'b010110100010101010: oled_data = 16'b1010101000101000;
				18'b010110100100101010: oled_data = 16'b1010101000001000;
				18'b010110100110101010: oled_data = 16'b1010101000001000;
				18'b010100011000101011: oled_data = 16'b1101110011010101;
				18'b010100011010101011: oled_data = 16'b1101110011010101;
				18'b010100011100101011: oled_data = 16'b1101110011010101;
				18'b010100011110101011: oled_data = 16'b1101110010110101;
				18'b010100100000101011: oled_data = 16'b1101010001110100;
				18'b010100100010101011: oled_data = 16'b1011001110010001;
				18'b010100100100101011: oled_data = 16'b1011001110010001;
				18'b010100100110101011: oled_data = 16'b1101010010010101;
				18'b010100101000101011: oled_data = 16'b1101010001010100;
				18'b010100101010101011: oled_data = 16'b1100110000010011;
				18'b010100101100101011: oled_data = 16'b1110010011010110;
				18'b010100101110101011: oled_data = 16'b1110010011010110;
				18'b010100110000101011: oled_data = 16'b1110010011010110;
				18'b010100110010101011: oled_data = 16'b1110010011010110;
				18'b010100110100101011: oled_data = 16'b1110010011010110;
				18'b010100110110101011: oled_data = 16'b1110010011110110;
				18'b010100111000101011: oled_data = 16'b1101010001110100;
				18'b010100111010101011: oled_data = 16'b1101110101110111;
				18'b010100111100101011: oled_data = 16'b1110111100011010;
				18'b010100111110101011: oled_data = 16'b1110111100011010;
				18'b010101000000101011: oled_data = 16'b1110111100011010;
				18'b010101000010101011: oled_data = 16'b1110111100011010;
				18'b010101000100101011: oled_data = 16'b1110111100011010;
				18'b010101000110101011: oled_data = 16'b1110011100011010;
				18'b010101001000101011: oled_data = 16'b1110011100011010;
				18'b010101001010101011: oled_data = 16'b1110111100011010;
				18'b010101001100101011: oled_data = 16'b1110111100011010;
				18'b010101001110101011: oled_data = 16'b1110111101011100;
				18'b010101010000101011: oled_data = 16'b1010010010110010;
				18'b010101010010101011: oled_data = 16'b0011000100100100;
				18'b010101010100101011: oled_data = 16'b0110001010101010;
				18'b010101010110101011: oled_data = 16'b1101111010111010;
				18'b010101011000101011: oled_data = 16'b1110111100111011;
				18'b010101011010101011: oled_data = 16'b1110111100011010;
				18'b010101011100101011: oled_data = 16'b1110111100011010;
				18'b010101011110101011: oled_data = 16'b1110111100011011;
				18'b010101100000101011: oled_data = 16'b1110111100011010;
				18'b010101100010101011: oled_data = 16'b1110111100011010;
				18'b010101100100101011: oled_data = 16'b1110111100011010;
				18'b010101100110101011: oled_data = 16'b1110111100011010;
				18'b010101101000101011: oled_data = 16'b1110111100011010;
				18'b010101101010101011: oled_data = 16'b1110111100011010;
				18'b010101101100101011: oled_data = 16'b1110111100011010;
				18'b010101101110101011: oled_data = 16'b1110111100011011;
				18'b010101110000101011: oled_data = 16'b1101011000110111;
				18'b010101110010101011: oled_data = 16'b1101011001111000;
				18'b010101110100101011: oled_data = 16'b1110111100011010;
				18'b010101110110101011: oled_data = 16'b1110111100011010;
				18'b010101111000101011: oled_data = 16'b1110111100011011;
				18'b010101111010101011: oled_data = 16'b1110011011011010;
				18'b010101111100101011: oled_data = 16'b1101010100110100;
				18'b010101111110101011: oled_data = 16'b1011101100001100;
				18'b010110000000101011: oled_data = 16'b1010101000101001;
				18'b010110000010101011: oled_data = 16'b1101110001110001;
				18'b010110000100101011: oled_data = 16'b1100101101101110;
				18'b010110000110101011: oled_data = 16'b1011001000101001;
				18'b010110001000101011: oled_data = 16'b1011101001001001;
				18'b010110001010101011: oled_data = 16'b1011001001001001;
				18'b010110001100101011: oled_data = 16'b1011001001001001;
				18'b010110001110101011: oled_data = 16'b1011001000101001;
				18'b010110010000101011: oled_data = 16'b1010101011001011;
				18'b010110010010101011: oled_data = 16'b1011111010111010;
				18'b010110010100101011: oled_data = 16'b1011111011111100;
				18'b010110010110101011: oled_data = 16'b1011111011111011;
				18'b010110011000101011: oled_data = 16'b1011111011111100;
				18'b010110011010101011: oled_data = 16'b1100011100111100;
				18'b010110011100101011: oled_data = 16'b1011110011010010;
				18'b010110011110101011: oled_data = 16'b1010101000001000;
				18'b010110100000101011: oled_data = 16'b1010101000101000;
				18'b010110100010101011: oled_data = 16'b1010101000001000;
				18'b010110100100101011: oled_data = 16'b1010101000001000;
				18'b010110100110101011: oled_data = 16'b1010101000001000;
				18'b010100011000101100: oled_data = 16'b1101110011010101;
				18'b010100011010101100: oled_data = 16'b1101110011010101;
				18'b010100011100101100: oled_data = 16'b1101110011010101;
				18'b010100011110101100: oled_data = 16'b1101010010010100;
				18'b010100100000101100: oled_data = 16'b1100001111110010;
				18'b010100100010101100: oled_data = 16'b1011001101110000;
				18'b010100100100101100: oled_data = 16'b1011101110010001;
				18'b010100100110101100: oled_data = 16'b1101110010110101;
				18'b010100101000101100: oled_data = 16'b1100110000110011;
				18'b010100101010101100: oled_data = 16'b1100110000010011;
				18'b010100101100101100: oled_data = 16'b1110010011010110;
				18'b010100101110101100: oled_data = 16'b1101110011010101;
				18'b010100110000101100: oled_data = 16'b1101110011010101;
				18'b010100110010101100: oled_data = 16'b1101110011010101;
				18'b010100110100101100: oled_data = 16'b1101110011010101;
				18'b010100110110101100: oled_data = 16'b1101110011010101;
				18'b010100111000101100: oled_data = 16'b1101010001110100;
				18'b010100111010101100: oled_data = 16'b1101110110110111;
				18'b010100111100101100: oled_data = 16'b1110111100011011;
				18'b010100111110101100: oled_data = 16'b1110111100011010;
				18'b010101000000101100: oled_data = 16'b1110111100011011;
				18'b010101000010101100: oled_data = 16'b1110111100011010;
				18'b010101000100101100: oled_data = 16'b1110111100011010;
				18'b010101000110101100: oled_data = 16'b1110011100011010;
				18'b010101001000101100: oled_data = 16'b1110011100011010;
				18'b010101001010101100: oled_data = 16'b1110111100011010;
				18'b010101001100101100: oled_data = 16'b1110111101011011;
				18'b010101001110101100: oled_data = 16'b1010110100110011;
				18'b010101010000101100: oled_data = 16'b0011100101100110;
				18'b010101010010101100: oled_data = 16'b0101001001101001;
				18'b010101010100101100: oled_data = 16'b1101011001011000;
				18'b010101010110101100: oled_data = 16'b1110111100011011;
				18'b010101011000101100: oled_data = 16'b1110011011111010;
				18'b010101011010101100: oled_data = 16'b1110011100011010;
				18'b010101011100101100: oled_data = 16'b1110011100011010;
				18'b010101011110101100: oled_data = 16'b1110011100011010;
				18'b010101100000101100: oled_data = 16'b1110011100011010;
				18'b010101100010101100: oled_data = 16'b1110011100011010;
				18'b010101100100101100: oled_data = 16'b1110011100011010;
				18'b010101100110101100: oled_data = 16'b1110011100011010;
				18'b010101101000101100: oled_data = 16'b1110111100011010;
				18'b010101101010101100: oled_data = 16'b1110111100111010;
				18'b010101101100101100: oled_data = 16'b1110111011111010;
				18'b010101101110101100: oled_data = 16'b1101010110110110;
				18'b010101110000101100: oled_data = 16'b1101010111010110;
				18'b010101110010101100: oled_data = 16'b1110111100011011;
				18'b010101110100101100: oled_data = 16'b1110111100011010;
				18'b010101110110101100: oled_data = 16'b1110111100011010;
				18'b010101111000101100: oled_data = 16'b1110111100011010;
				18'b010101111010101100: oled_data = 16'b1110011100011010;
				18'b010101111100101100: oled_data = 16'b1101110101110101;
				18'b010101111110101100: oled_data = 16'b1011101011101100;
				18'b010110000000101100: oled_data = 16'b1011001001001010;
				18'b010110000010101100: oled_data = 16'b1101110010010010;
				18'b010110000100101100: oled_data = 16'b1100001011101100;
				18'b010110000110101100: oled_data = 16'b1011001000101001;
				18'b010110001000101100: oled_data = 16'b1011001001001001;
				18'b010110001010101100: oled_data = 16'b1011001001001001;
				18'b010110001100101100: oled_data = 16'b1011001001001001;
				18'b010110001110101100: oled_data = 16'b1011001000101001;
				18'b010110010000101100: oled_data = 16'b1011110000110001;
				18'b010110010010101100: oled_data = 16'b1100011100011100;
				18'b010110010100101100: oled_data = 16'b1011111011111011;
				18'b010110010110101100: oled_data = 16'b1011111011111011;
				18'b010110011000101100: oled_data = 16'b1011111011111100;
				18'b010110011010101100: oled_data = 16'b1100111100111101;
				18'b010110011100101100: oled_data = 16'b1011111000111000;
				18'b010110011110101100: oled_data = 16'b1010101010001010;
				18'b010110100000101100: oled_data = 16'b1010101000101000;
				18'b010110100010101100: oled_data = 16'b1010101000001000;
				18'b010110100100101100: oled_data = 16'b1010101000001000;
				18'b010110100110101100: oled_data = 16'b1010101000001000;
				18'b010100011000101101: oled_data = 16'b1101110010110101;
				18'b010100011010101101: oled_data = 16'b1101110010110101;
				18'b010100011100101101: oled_data = 16'b1101110010110101;
				18'b010100011110101101: oled_data = 16'b1100110001010011;
				18'b010100100000101101: oled_data = 16'b1011101110110001;
				18'b010100100010101101: oled_data = 16'b1011001101110000;
				18'b010100100100101101: oled_data = 16'b1011001110010001;
				18'b010100100110101101: oled_data = 16'b1101110010110101;
				18'b010100101000101101: oled_data = 16'b1100110000110011;
				18'b010100101010101101: oled_data = 16'b1100110000110011;
				18'b010100101100101101: oled_data = 16'b1101110011010110;
				18'b010100101110101101: oled_data = 16'b1101110010110101;
				18'b010100110000101101: oled_data = 16'b1101110010110101;
				18'b010100110010101101: oled_data = 16'b1101110010110101;
				18'b010100110100101101: oled_data = 16'b1101110010110101;
				18'b010100110110101101: oled_data = 16'b1101110010110101;
				18'b010100111000101101: oled_data = 16'b1100110001010011;
				18'b010100111010101101: oled_data = 16'b1101110111111000;
				18'b010100111100101101: oled_data = 16'b1110111100111011;
				18'b010100111110101101: oled_data = 16'b1110111100011010;
				18'b010101000000101101: oled_data = 16'b1110111100011010;
				18'b010101000010101101: oled_data = 16'b1110111100011010;
				18'b010101000100101101: oled_data = 16'b1110111100011010;
				18'b010101000110101101: oled_data = 16'b1110111100011010;
				18'b010101001000101101: oled_data = 16'b1110111100011010;
				18'b010101001010101101: oled_data = 16'b1110111100111010;
				18'b010101001100101101: oled_data = 16'b1100010111010101;
				18'b010101001110101101: oled_data = 16'b0100000110100110;
				18'b010101010000101101: oled_data = 16'b0100101000101000;
				18'b010101010010101101: oled_data = 16'b1100011000010111;
				18'b010101010100101101: oled_data = 16'b1110111100111011;
				18'b010101010110101101: oled_data = 16'b1110011011111010;
				18'b010101011000101101: oled_data = 16'b1110111011111010;
				18'b010101011010101101: oled_data = 16'b1110111011111010;
				18'b010101011100101101: oled_data = 16'b1110011100011010;
				18'b010101011110101101: oled_data = 16'b1110011100011010;
				18'b010101100000101101: oled_data = 16'b1110011100011010;
				18'b010101100010101101: oled_data = 16'b1110011100011010;
				18'b010101100100101101: oled_data = 16'b1110011100011010;
				18'b010101100110101101: oled_data = 16'b1110111100011010;
				18'b010101101000101101: oled_data = 16'b1110111100011010;
				18'b010101101010101101: oled_data = 16'b1101111000010111;
				18'b010101101100101101: oled_data = 16'b1101010101010101;
				18'b010101101110101101: oled_data = 16'b1101110101010101;
				18'b010101110000101101: oled_data = 16'b1110111011011010;
				18'b010101110010101101: oled_data = 16'b1110111100011011;
				18'b010101110100101101: oled_data = 16'b1110111100011010;
				18'b010101110110101101: oled_data = 16'b1110111100011010;
				18'b010101111000101101: oled_data = 16'b1110111100011010;
				18'b010101111010101101: oled_data = 16'b1110111100011010;
				18'b010101111100101101: oled_data = 16'b1101010110010110;
				18'b010101111110101101: oled_data = 16'b1011101011001100;
				18'b010110000000101101: oled_data = 16'b1011001001001010;
				18'b010110000010101101: oled_data = 16'b1101110001010001;
				18'b010110000100101101: oled_data = 16'b1011101010101011;
				18'b010110000110101101: oled_data = 16'b1011001001001001;
				18'b010110001000101101: oled_data = 16'b1011001001001001;
				18'b010110001010101101: oled_data = 16'b1011001001001001;
				18'b010110001100101101: oled_data = 16'b1011001001001001;
				18'b010110001110101101: oled_data = 16'b1011001001001001;
				18'b010110010000101101: oled_data = 16'b1100010110010111;
				18'b010110010010101101: oled_data = 16'b1011111100011100;
				18'b010110010100101101: oled_data = 16'b1011111011111011;
				18'b010110010110101101: oled_data = 16'b1011111011111011;
				18'b010110011000101101: oled_data = 16'b1011111011111100;
				18'b010110011010101101: oled_data = 16'b1100111100011101;
				18'b010110011100101101: oled_data = 16'b1011111011111011;
				18'b010110011110101101: oled_data = 16'b1010101101101101;
				18'b010110100000101101: oled_data = 16'b1010101000001000;
				18'b010110100010101101: oled_data = 16'b1010101000001000;
				18'b010110100100101101: oled_data = 16'b1010101000001000;
				18'b010110100110101101: oled_data = 16'b1010101000001000;
				18'b010100011000101110: oled_data = 16'b1101110010110101;
				18'b010100011010101110: oled_data = 16'b1101110010110101;
				18'b010100011100101110: oled_data = 16'b1101110010110101;
				18'b010100011110101110: oled_data = 16'b1100110000010011;
				18'b010100100000101110: oled_data = 16'b1011001110010001;
				18'b010100100010101110: oled_data = 16'b1011001101010000;
				18'b010100100100101110: oled_data = 16'b1011101110110001;
				18'b010100100110101110: oled_data = 16'b1101110010110101;
				18'b010100101000101110: oled_data = 16'b1100001111110010;
				18'b010100101010101110: oled_data = 16'b1100110000110011;
				18'b010100101100101110: oled_data = 16'b1101110011010110;
				18'b010100101110101110: oled_data = 16'b1101110010110101;
				18'b010100110000101110: oled_data = 16'b1101110010110101;
				18'b010100110010101110: oled_data = 16'b1101110010110101;
				18'b010100110100101110: oled_data = 16'b1101110010110101;
				18'b010100110110101110: oled_data = 16'b1101110010110101;
				18'b010100111000101110: oled_data = 16'b1100110001110011;
				18'b010100111010101110: oled_data = 16'b1101111000111000;
				18'b010100111100101110: oled_data = 16'b1110011100011010;
				18'b010100111110101110: oled_data = 16'b1110011100011010;
				18'b010101000000101110: oled_data = 16'b1110011011111010;
				18'b010101000010101110: oled_data = 16'b1110011011111010;
				18'b010101000100101110: oled_data = 16'b1110011100011010;
				18'b010101000110101110: oled_data = 16'b1110011100011010;
				18'b010101001000101110: oled_data = 16'b1110011100011010;
				18'b010101001010101110: oled_data = 16'b1101111011011001;
				18'b010101001100101110: oled_data = 16'b1100110111110110;
				18'b010101001110101110: oled_data = 16'b1010010011010001;
				18'b010101010000101110: oled_data = 16'b1101011001011000;
				18'b010101010010101110: oled_data = 16'b1110111100111011;
				18'b010101010100101110: oled_data = 16'b1110111100011010;
				18'b010101010110101110: oled_data = 16'b1110111100011010;
				18'b010101011000101110: oled_data = 16'b1110111100011010;
				18'b010101011010101110: oled_data = 16'b1110111100011010;
				18'b010101011100101110: oled_data = 16'b1110011100011010;
				18'b010101011110101110: oled_data = 16'b1110011100011010;
				18'b010101100000101110: oled_data = 16'b1110011100011010;
				18'b010101100010101110: oled_data = 16'b1110111100011010;
				18'b010101100100101110: oled_data = 16'b1110111100011010;
				18'b010101100110101110: oled_data = 16'b1101111001011000;
				18'b010101101000101110: oled_data = 16'b1100010011110011;
				18'b010101101010101110: oled_data = 16'b1100110010010010;
				18'b010101101100101110: oled_data = 16'b1101110100010100;
				18'b010101101110101110: oled_data = 16'b1110011000111000;
				18'b010101110000101110: oled_data = 16'b1110111100011010;
				18'b010101110010101110: oled_data = 16'b1110111100011010;
				18'b010101110100101110: oled_data = 16'b1110111100011010;
				18'b010101110110101110: oled_data = 16'b1110111100011010;
				18'b010101111000101110: oled_data = 16'b1110011100011010;
				18'b010101111010101110: oled_data = 16'b1110011100011010;
				18'b010101111100101110: oled_data = 16'b1101111000110111;
				18'b010101111110101110: oled_data = 16'b1011001011001011;
				18'b010110000000101110: oled_data = 16'b1011001001101010;
				18'b010110000010101110: oled_data = 16'b1101010000110000;
				18'b010110000100101110: oled_data = 16'b1011101001101010;
				18'b010110000110101110: oled_data = 16'b1011001001001001;
				18'b010110001000101110: oled_data = 16'b1011001000101001;
				18'b010110001010101110: oled_data = 16'b1011001001001001;
				18'b010110001100101110: oled_data = 16'b1011001000101001;
				18'b010110001110101110: oled_data = 16'b1011001010001010;
				18'b010110010000101110: oled_data = 16'b1100011001011001;
				18'b010110010010101110: oled_data = 16'b1011111011111100;
				18'b010110010100101110: oled_data = 16'b1011111011011011;
				18'b010110010110101110: oled_data = 16'b1011111011011011;
				18'b010110011000101110: oled_data = 16'b1011111011011011;
				18'b010110011010101110: oled_data = 16'b1100111100011100;
				18'b010110011100101110: oled_data = 16'b1011111100011100;
				18'b010110011110101110: oled_data = 16'b1011010010010010;
				18'b010110100000101110: oled_data = 16'b1010100111101000;
				18'b010110100010101110: oled_data = 16'b1010101000001000;
				18'b010110100100101110: oled_data = 16'b1010101000001000;
				18'b010110100110101110: oled_data = 16'b1010101000001000;
				18'b010100011000101111: oled_data = 16'b1101110010010101;
				18'b010100011010101111: oled_data = 16'b1101110010010101;
				18'b010100011100101111: oled_data = 16'b1101010010010101;
				18'b010100011110101111: oled_data = 16'b1100001111010010;
				18'b010100100000101111: oled_data = 16'b1011001101010000;
				18'b010100100010101111: oled_data = 16'b1011001101010000;
				18'b010100100100101111: oled_data = 16'b1011101111010010;
				18'b010100100110101111: oled_data = 16'b1101110011010101;
				18'b010100101000101111: oled_data = 16'b1011101111010001;
				18'b010100101010101111: oled_data = 16'b1100110000010010;
				18'b010100101100101111: oled_data = 16'b1101110011010110;
				18'b010100101110101111: oled_data = 16'b1101110010110101;
				18'b010100110000101111: oled_data = 16'b1101110010110101;
				18'b010100110010101111: oled_data = 16'b1101110010110101;
				18'b010100110100101111: oled_data = 16'b1101110010110101;
				18'b010100110110101111: oled_data = 16'b1101110010110101;
				18'b010100111000101111: oled_data = 16'b1100110001110011;
				18'b010100111010101111: oled_data = 16'b1101111001111001;
				18'b010100111100101111: oled_data = 16'b1110011100111010;
				18'b010100111110101111: oled_data = 16'b1110011011111010;
				18'b010101000000101111: oled_data = 16'b1110011100011010;
				18'b010101000010101111: oled_data = 16'b1110011100011010;
				18'b010101000100101111: oled_data = 16'b1110011100011010;
				18'b010101000110101111: oled_data = 16'b1110011011111010;
				18'b010101001000101111: oled_data = 16'b1110011011111010;
				18'b010101001010101111: oled_data = 16'b1110011011111010;
				18'b010101001100101111: oled_data = 16'b1110111100011010;
				18'b010101001110101111: oled_data = 16'b1110111100111011;
				18'b010101010000101111: oled_data = 16'b1110111100011010;
				18'b010101010010101111: oled_data = 16'b1110011100011010;
				18'b010101010100101111: oled_data = 16'b1110011100011010;
				18'b010101010110101111: oled_data = 16'b1110011100011010;
				18'b010101011000101111: oled_data = 16'b1110011100011010;
				18'b010101011010101111: oled_data = 16'b1110111100011010;
				18'b010101011100101111: oled_data = 16'b1110111100011010;
				18'b010101011110101111: oled_data = 16'b1110111100011010;
				18'b010101100000101111: oled_data = 16'b1110011011011001;
				18'b010101100010101111: oled_data = 16'b1101010111010110;
				18'b010101100100101111: oled_data = 16'b1011110010110010;
				18'b010101100110101111: oled_data = 16'b1011001111001111;
				18'b010101101000101111: oled_data = 16'b1100010000110001;
				18'b010101101010101111: oled_data = 16'b1101110100010101;
				18'b010101101100101111: oled_data = 16'b1101010100010100;
				18'b010101101110101111: oled_data = 16'b1110011010011001;
				18'b010101110000101111: oled_data = 16'b1110011011111010;
				18'b010101110010101111: oled_data = 16'b1110011011111010;
				18'b010101110100101111: oled_data = 16'b1110011011111010;
				18'b010101110110101111: oled_data = 16'b1110011011111010;
				18'b010101111000101111: oled_data = 16'b1110011011111010;
				18'b010101111010101111: oled_data = 16'b1110011100011010;
				18'b010101111100101111: oled_data = 16'b1110011011111001;
				18'b010101111110101111: oled_data = 16'b1010101100101100;
				18'b010110000000101111: oled_data = 16'b1011001001101010;
				18'b010110000010101111: oled_data = 16'b1100101111101111;
				18'b010110000100101111: oled_data = 16'b1011001001001001;
				18'b010110000110101111: oled_data = 16'b1011001000101001;
				18'b010110001000101111: oled_data = 16'b1011001001101001;
				18'b010110001010101111: oled_data = 16'b1011001001001001;
				18'b010110001100101111: oled_data = 16'b1011001000101000;
				18'b010110001110101111: oled_data = 16'b1011101011101100;
				18'b010110010000101111: oled_data = 16'b1100011010111011;
				18'b010110010010101111: oled_data = 16'b1011111011011100;
				18'b010110010100101111: oled_data = 16'b1011111011011011;
				18'b010110010110101111: oled_data = 16'b1011111011011011;
				18'b010110011000101111: oled_data = 16'b1011111011011100;
				18'b010110011010101111: oled_data = 16'b1100011011111100;
				18'b010110011100101111: oled_data = 16'b1011111100011100;
				18'b010110011110101111: oled_data = 16'b1011110100010100;
				18'b010110100000101111: oled_data = 16'b1010100111101000;
				18'b010110100010101111: oled_data = 16'b1010100111101000;
				18'b010110100100101111: oled_data = 16'b1010101000001000;
				18'b010110100110101111: oled_data = 16'b1010100111101000;
				18'b010100011000110000: oled_data = 16'b1101010001110100;
				18'b010100011010110000: oled_data = 16'b1101010001110100;
				18'b010100011100110000: oled_data = 16'b1101010001010100;
				18'b010100011110110000: oled_data = 16'b1011101110010001;
				18'b010100100000110000: oled_data = 16'b1010101100101111;
				18'b010100100010110000: oled_data = 16'b1010101100101111;
				18'b010100100100110000: oled_data = 16'b1011101111010010;
				18'b010100100110110000: oled_data = 16'b1101110010110101;
				18'b010100101000110000: oled_data = 16'b1011101110110001;
				18'b010100101010110000: oled_data = 16'b1100010000010010;
				18'b010100101100110000: oled_data = 16'b1101110011010101;
				18'b010100101110110000: oled_data = 16'b1101110010110101;
				18'b010100110000110000: oled_data = 16'b1101010001110100;
				18'b010100110010110000: oled_data = 16'b1101010010010100;
				18'b010100110100110000: oled_data = 16'b1101110010110101;
				18'b010100110110110000: oled_data = 16'b1101110010110101;
				18'b010100111000110000: oled_data = 16'b1100110010010100;
				18'b010100111010110000: oled_data = 16'b1110011001111001;
				18'b010100111100110000: oled_data = 16'b1100110101110101;
				18'b010100111110110000: oled_data = 16'b1010110001010001;
				18'b010101000000110000: oled_data = 16'b1100110101110101;
				18'b010101000010110000: oled_data = 16'b1101111001111000;
				18'b010101000100110000: oled_data = 16'b1110011011111010;
				18'b010101000110110000: oled_data = 16'b1110011100011010;
				18'b010101001000110000: oled_data = 16'b1110011011111010;
				18'b010101001010110000: oled_data = 16'b1110011011111010;
				18'b010101001100110000: oled_data = 16'b1110011011111010;
				18'b010101001110110000: oled_data = 16'b1110011011111010;
				18'b010101010000110000: oled_data = 16'b1110011100011010;
				18'b010101010010110000: oled_data = 16'b1110011100011010;
				18'b010101010100110000: oled_data = 16'b1110111100011010;
				18'b010101010110110000: oled_data = 16'b1110111100011010;
				18'b010101011000110000: oled_data = 16'b1110011011111010;
				18'b010101011010110000: oled_data = 16'b1101111001111000;
				18'b010101011100110000: oled_data = 16'b1101010111010110;
				18'b010101011110110000: oled_data = 16'b1100010100010100;
				18'b010101100000110000: oled_data = 16'b1011110000110001;
				18'b010101100010110000: oled_data = 16'b1011001110101111;
				18'b010101100100110000: oled_data = 16'b1011101110110000;
				18'b010101100110110000: oled_data = 16'b1100110001010010;
				18'b010101101000110000: oled_data = 16'b1101110100010100;
				18'b010101101010110000: oled_data = 16'b1101010010110011;
				18'b010101101100110000: oled_data = 16'b1101010011110100;
				18'b010101101110110000: oled_data = 16'b1100110110010101;
				18'b010101110000110000: oled_data = 16'b1101111010111001;
				18'b010101110010110000: oled_data = 16'b1110011011111010;
				18'b010101110100110000: oled_data = 16'b1110011011111010;
				18'b010101110110110000: oled_data = 16'b1110011011111010;
				18'b010101111000110000: oled_data = 16'b1110011011111010;
				18'b010101111010110000: oled_data = 16'b1110011011111010;
				18'b010101111100110000: oled_data = 16'b1110011011111010;
				18'b010101111110110000: oled_data = 16'b1011001110101110;
				18'b010110000000110000: oled_data = 16'b1011001001101010;
				18'b010110000010110000: oled_data = 16'b1100101110001110;
				18'b010110000100110000: oled_data = 16'b1011001000101001;
				18'b010110000110110000: oled_data = 16'b1011001000101001;
				18'b010110001000110000: oled_data = 16'b1100101101101101;
				18'b010110001010110000: oled_data = 16'b1011101001101010;
				18'b010110001100110000: oled_data = 16'b1011001000101000;
				18'b010110001110110000: oled_data = 16'b1011101100001100;
				18'b010110010000110000: oled_data = 16'b1100011010111011;
				18'b010110010010110000: oled_data = 16'b1011111011011100;
				18'b010110010100110000: oled_data = 16'b1011111011011100;
				18'b010110010110110000: oled_data = 16'b1011011010111011;
				18'b010110011000110000: oled_data = 16'b1010111001111010;
				18'b010110011010110000: oled_data = 16'b1011011010111011;
				18'b010110011100110000: oled_data = 16'b1011111100011100;
				18'b010110011110110000: oled_data = 16'b1011110100110101;
				18'b010110100000110000: oled_data = 16'b1010100111001000;
				18'b010110100010110000: oled_data = 16'b1001100111000111;
				18'b010110100100110000: oled_data = 16'b1001100111000111;
				18'b010110100110110000: oled_data = 16'b1001100111000111;
				18'b010100011000110001: oled_data = 16'b1101010001010100;
				18'b010100011010110001: oled_data = 16'b1101010001010100;
				18'b010100011100110001: oled_data = 16'b1100001111110010;
				18'b010100011110110001: oled_data = 16'b1010101100101111;
				18'b010100100000110001: oled_data = 16'b1010101100001111;
				18'b010100100010110001: oled_data = 16'b1010101100001111;
				18'b010100100100110001: oled_data = 16'b1100001111010010;
				18'b010100100110110001: oled_data = 16'b1101110010110101;
				18'b010100101000110001: oled_data = 16'b1011101110110001;
				18'b010100101010110001: oled_data = 16'b1100001111110010;
				18'b010100101100110001: oled_data = 16'b1101110010110101;
				18'b010100101110110001: oled_data = 16'b1101010010010100;
				18'b010100110000110001: oled_data = 16'b1101010001010100;
				18'b010100110010110001: oled_data = 16'b1100110000110100;
				18'b010100110100110001: oled_data = 16'b1101010010010101;
				18'b010100110110110001: oled_data = 16'b1101110010010101;
				18'b010100111000110001: oled_data = 16'b1100110001010100;
				18'b010100111010110001: oled_data = 16'b1011010000010001;
				18'b010100111100110001: oled_data = 16'b1011001101101111;
				18'b010100111110110001: oled_data = 16'b1011001101110000;
				18'b010101000000110001: oled_data = 16'b1010101101001111;
				18'b010101000010110001: oled_data = 16'b1011001110110000;
				18'b010101000100110001: oled_data = 16'b1011110000110001;
				18'b010101000110110001: oled_data = 16'b1011110011010011;
				18'b010101001000110001: oled_data = 16'b1100010101110101;
				18'b010101001010110001: oled_data = 16'b1100111000110111;
				18'b010101001100110001: oled_data = 16'b1101011001010111;
				18'b010101001110110001: oled_data = 16'b1100111000110111;
				18'b010101010000110001: oled_data = 16'b1011110110110101;
				18'b010101010010110001: oled_data = 16'b1100110101110101;
				18'b010101010100110001: oled_data = 16'b1100010100110100;
				18'b010101010110110001: oled_data = 16'b1011110010110010;
				18'b010101011000110001: oled_data = 16'b1011010000110001;
				18'b010101011010110001: oled_data = 16'b1010101110101111;
				18'b010101011100110001: oled_data = 16'b1011001110001111;
				18'b010101011110110001: oled_data = 16'b1011101110101111;
				18'b010101100000110001: oled_data = 16'b1011101110110000;
				18'b010101100010110001: oled_data = 16'b1011101111010000;
				18'b010101100100110001: oled_data = 16'b1100110001110010;
				18'b010101100110110001: oled_data = 16'b1101110100010101;
				18'b010101101000110001: oled_data = 16'b1101010011010100;
				18'b010101101010110001: oled_data = 16'b1101010011010100;
				18'b010101101100110001: oled_data = 16'b1100110010110011;
				18'b010101101110110001: oled_data = 16'b1100110100110100;
				18'b010101110000110001: oled_data = 16'b1101111001111001;
				18'b010101110010110001: oled_data = 16'b1110011011111010;
				18'b010101110100110001: oled_data = 16'b1110011011011010;
				18'b010101110110110001: oled_data = 16'b1110011011011010;
				18'b010101111000110001: oled_data = 16'b1110011011111010;
				18'b010101111010110001: oled_data = 16'b1110011011011001;
				18'b010101111100110001: oled_data = 16'b1110011011011001;
				18'b010101111110110001: oled_data = 16'b1011001111001110;
				18'b010110000000110001: oled_data = 16'b1011001001101001;
				18'b010110000010110001: oled_data = 16'b1100001101001101;
				18'b010110000100110001: oled_data = 16'b1011001000101001;
				18'b010110000110110001: oled_data = 16'b1011001001001001;
				18'b010110001000110001: oled_data = 16'b1100101101101101;
				18'b010110001010110001: oled_data = 16'b1011001001001001;
				18'b010110001100110001: oled_data = 16'b1011001000001000;
				18'b010110001110110001: oled_data = 16'b1011101011101100;
				18'b010110010000110001: oled_data = 16'b1100011010111011;
				18'b010110010010110001: oled_data = 16'b1011111011111100;
				18'b010110010100110001: oled_data = 16'b1011011011011011;
				18'b010110010110110001: oled_data = 16'b1001110111111000;
				18'b010110011000110001: oled_data = 16'b1001010110111000;
				18'b010110011010110001: oled_data = 16'b1010111001111010;
				18'b010110011100110001: oled_data = 16'b1011111100011100;
				18'b010110011110110001: oled_data = 16'b1011010010010010;
				18'b010110100000110001: oled_data = 16'b1010000111000111;
				18'b010110100010110001: oled_data = 16'b1010100111101000;
				18'b010110100100110001: oled_data = 16'b1010000111100111;
				18'b010110100110110001: oled_data = 16'b1010000111000111;
				18'b010100011000110010: oled_data = 16'b1100110001010100;
				18'b010100011010110010: oled_data = 16'b1101010001010100;
				18'b010100011100110010: oled_data = 16'b1011101111010010;
				18'b010100011110110010: oled_data = 16'b1010101100001111;
				18'b010100100000110010: oled_data = 16'b1010001100001111;
				18'b010100100010110010: oled_data = 16'b1010001011101110;
				18'b010100100100110010: oled_data = 16'b1011101111010010;
				18'b010100100110110010: oled_data = 16'b1101010001110100;
				18'b010100101000110010: oled_data = 16'b1011101110010001;
				18'b010100101010110010: oled_data = 16'b1011101110110001;
				18'b010100101100110010: oled_data = 16'b1101010010010101;
				18'b010100101110110010: oled_data = 16'b1101010001110100;
				18'b010100110000110010: oled_data = 16'b1101010001010100;
				18'b010100110010110010: oled_data = 16'b1100110000010011;
				18'b010100110100110010: oled_data = 16'b1101010001110100;
				18'b010100110110110010: oled_data = 16'b1101010001110100;
				18'b010100111000110010: oled_data = 16'b1011101111010001;
				18'b010100111010110010: oled_data = 16'b1010101101001111;
				18'b010100111100110010: oled_data = 16'b1011101110010000;
				18'b010100111110110010: oled_data = 16'b1011001110010000;
				18'b010101000000110010: oled_data = 16'b1011001101110000;
				18'b010101000010110010: oled_data = 16'b1011001101101111;
				18'b010101000100110010: oled_data = 16'b1010101101001110;
				18'b010101000110110010: oled_data = 16'b1011110000110001;
				18'b010101001000110010: oled_data = 16'b1101110111110111;
				18'b010101001010110010: oled_data = 16'b1101111010011001;
				18'b010101001100110010: oled_data = 16'b1101111010111001;
				18'b010101001110110010: oled_data = 16'b1101111010011000;
				18'b010101010000110010: oled_data = 16'b1100110111010110;
				18'b010101010010110010: oled_data = 16'b1011110001110010;
				18'b010101010100110010: oled_data = 16'b1011001111010000;
				18'b010101010110110010: oled_data = 16'b1011001110001111;
				18'b010101011000110010: oled_data = 16'b1011001110001111;
				18'b010101011010110010: oled_data = 16'b1011001110001111;
				18'b010101011100110010: oled_data = 16'b1011101110101111;
				18'b010101011110110010: oled_data = 16'b1011101110110000;
				18'b010101100000110010: oled_data = 16'b1100010000010001;
				18'b010101100010110010: oled_data = 16'b1100010000110001;
				18'b010101100100110010: oled_data = 16'b1101110011010100;
				18'b010101100110110010: oled_data = 16'b1101010010110011;
				18'b010101101000110010: oled_data = 16'b1100110010010011;
				18'b010101101010110010: oled_data = 16'b1101110011110101;
				18'b010101101100110010: oled_data = 16'b1100110010010011;
				18'b010101101110110010: oled_data = 16'b1100010011010011;
				18'b010101110000110010: oled_data = 16'b1101010111010111;
				18'b010101110010110010: oled_data = 16'b1110011010011001;
				18'b010101110100110010: oled_data = 16'b1110011010111001;
				18'b010101110110110010: oled_data = 16'b1110011010111001;
				18'b010101111000110010: oled_data = 16'b1101111001111000;
				18'b010101111010110010: oled_data = 16'b1101011001011000;
				18'b010101111100110010: oled_data = 16'b1110011001111000;
				18'b010101111110110010: oled_data = 16'b1011001110001101;
				18'b010110000000110010: oled_data = 16'b1011001001001001;
				18'b010110000010110010: oled_data = 16'b1100001100101100;
				18'b010110000100110010: oled_data = 16'b1011001000101001;
				18'b010110000110110010: oled_data = 16'b1011001001001001;
				18'b010110001000110010: oled_data = 16'b1011101010101010;
				18'b010110001010110010: oled_data = 16'b1011001000101000;
				18'b010110001100110010: oled_data = 16'b1011001000001000;
				18'b010110001110110010: oled_data = 16'b1011001001101010;
				18'b010110010000110010: oled_data = 16'b1100011001011001;
				18'b010110010010110010: oled_data = 16'b1011111011111100;
				18'b010110010100110010: oled_data = 16'b1010011000111001;
				18'b010110010110110010: oled_data = 16'b1001010110110111;
				18'b010110011000110010: oled_data = 16'b1000110110110111;
				18'b010110011010110010: oled_data = 16'b1001110111111000;
				18'b010110011100110010: oled_data = 16'b1010111010011010;
				18'b010110011110110010: oled_data = 16'b1010101110101110;
				18'b010110100000110010: oled_data = 16'b1010000110100111;
				18'b010110100010110010: oled_data = 16'b1010000111000111;
				18'b010110100100110010: oled_data = 16'b1010000111000111;
				18'b010110100110110010: oled_data = 16'b1010000111000111;
				18'b010100011000110011: oled_data = 16'b1100110000110011;
				18'b010100011010110011: oled_data = 16'b1100110000110011;
				18'b010100011100110011: oled_data = 16'b1011001101010000;
				18'b010100011110110011: oled_data = 16'b1010001011101110;
				18'b010100100000110011: oled_data = 16'b1010001011101110;
				18'b010100100010110011: oled_data = 16'b1010001011001110;
				18'b010100100100110011: oled_data = 16'b1011001110010001;
				18'b010100100110110011: oled_data = 16'b1100110001010100;
				18'b010100101000110011: oled_data = 16'b1011001110010001;
				18'b010100101010110011: oled_data = 16'b1011001101010000;
				18'b010100101100110011: oled_data = 16'b1100110001010100;
				18'b010100101110110011: oled_data = 16'b1100110001010100;
				18'b010100110000110011: oled_data = 16'b1100110000110100;
				18'b010100110010110011: oled_data = 16'b1100001111110010;
				18'b010100110100110011: oled_data = 16'b1100110001010100;
				18'b010100110110110011: oled_data = 16'b1101010001010100;
				18'b010100111000110011: oled_data = 16'b1011001110010000;
				18'b010100111010110011: oled_data = 16'b1010001011101110;
				18'b010100111100110011: oled_data = 16'b1010101100101110;
				18'b010100111110110011: oled_data = 16'b1010101101001111;
				18'b010101000000110011: oled_data = 16'b1010101101101111;
				18'b010101000010110011: oled_data = 16'b1010101101001110;
				18'b010101000100110011: oled_data = 16'b1011010001110001;
				18'b010101000110110011: oled_data = 16'b1101111010011001;
				18'b010101001000110011: oled_data = 16'b1101111010111001;
				18'b010101001010110011: oled_data = 16'b1101111010111001;
				18'b010101001100110011: oled_data = 16'b1110011010011001;
				18'b010101001110110011: oled_data = 16'b1101111010111001;
				18'b010101010000110011: oled_data = 16'b1110011010111001;
				18'b010101010010110011: oled_data = 16'b1101111001011000;
				18'b010101010100110011: oled_data = 16'b1011110100010011;
				18'b010101010110110011: oled_data = 16'b1010101111001111;
				18'b010101011000110011: oled_data = 16'b1011001110001111;
				18'b010101011010110011: oled_data = 16'b1011001110001111;
				18'b010101011100110011: oled_data = 16'b1011101111010000;
				18'b010101011110110011: oled_data = 16'b1100110001110010;
				18'b010101100000110011: oled_data = 16'b1101010010110011;
				18'b010101100010110011: oled_data = 16'b1100010000110010;
				18'b010101100100110011: oled_data = 16'b1100110010010010;
				18'b010101100110110011: oled_data = 16'b1100110010010011;
				18'b010101101000110011: oled_data = 16'b1101010011110100;
				18'b010101101010110011: oled_data = 16'b1101010011010101;
				18'b010101101100110011: oled_data = 16'b1100110010110011;
				18'b010101101110110011: oled_data = 16'b1100110010010011;
				18'b010101110000110011: oled_data = 16'b1100110011110100;
				18'b010101110010110011: oled_data = 16'b1100110101010101;
				18'b010101110100110011: oled_data = 16'b1100110110110110;
				18'b010101110110110011: oled_data = 16'b1100110111110110;
				18'b010101111000110011: oled_data = 16'b1101010111110111;
				18'b010101111010110011: oled_data = 16'b1101110110110111;
				18'b010101111100110011: oled_data = 16'b1101010100110100;
				18'b010101111110110011: oled_data = 16'b1011001100001100;
				18'b010110000000110011: oled_data = 16'b1011001000101001;
				18'b010110000010110011: oled_data = 16'b1011101100001100;
				18'b010110000100110011: oled_data = 16'b1010101000001000;
				18'b010110000110110011: oled_data = 16'b1011001000001000;
				18'b010110001000110011: oled_data = 16'b1011001000001000;
				18'b010110001010110011: oled_data = 16'b1011001000001000;
				18'b010110001100110011: oled_data = 16'b1010101000001000;
				18'b010110001110110011: oled_data = 16'b1011001000001000;
				18'b010110010000110011: oled_data = 16'b1011110100010100;
				18'b010110010010110011: oled_data = 16'b1011011011111011;
				18'b010110010100110011: oled_data = 16'b1001010111010111;
				18'b010110010110110011: oled_data = 16'b1000110110010110;
				18'b010110011000110011: oled_data = 16'b1000110110010111;
				18'b010110011010110011: oled_data = 16'b1000110101110111;
				18'b010110011100110011: oled_data = 16'b1010010111010111;
				18'b010110011110110011: oled_data = 16'b1010001001101010;
				18'b010110100000110011: oled_data = 16'b1010000111000111;
				18'b010110100010110011: oled_data = 16'b1001100111000111;
				18'b010110100100110011: oled_data = 16'b1001100111000111;
				18'b010110100110110011: oled_data = 16'b1001100111000111;
				18'b010100011000110100: oled_data = 16'b1100110000010011;
				18'b010100011010110100: oled_data = 16'b1100110000010011;
				18'b010100011100110100: oled_data = 16'b1010101011101111;
				18'b010100011110110100: oled_data = 16'b1001101010101101;
				18'b010100100000110100: oled_data = 16'b1001101010101110;
				18'b010100100010110100: oled_data = 16'b1001101011001110;
				18'b010100100100110100: oled_data = 16'b1011001110010000;
				18'b010100100110110100: oled_data = 16'b1100110000110011;
				18'b010100101000110100: oled_data = 16'b1011001101110000;
				18'b010100101010110100: oled_data = 16'b1010001011101111;
				18'b010100101100110100: oled_data = 16'b1100110000010011;
				18'b010100101110110100: oled_data = 16'b1100110000010011;
				18'b010100110000110100: oled_data = 16'b1100110000010011;
				18'b010100110010110100: oled_data = 16'b1100001111010010;
				18'b010100110100110100: oled_data = 16'b1100110000110011;
				18'b010100110110110100: oled_data = 16'b1100110000110011;
				18'b010100111000110100: oled_data = 16'b1011001110010000;
				18'b010100111010110100: oled_data = 16'b1010001100001110;
				18'b010100111100110100: oled_data = 16'b1010101100101110;
				18'b010100111110110100: oled_data = 16'b1010001100001110;
				18'b010101000000110100: oled_data = 16'b1010001011101101;
				18'b010101000010110100: oled_data = 16'b1010101110101111;
				18'b010101000100110100: oled_data = 16'b1101111001011000;
				18'b010101000110110100: oled_data = 16'b1101111010111001;
				18'b010101001000110100: oled_data = 16'b1101111010111001;
				18'b010101001010110100: oled_data = 16'b1101111010011001;
				18'b010101001100110100: oled_data = 16'b1110011010011001;
				18'b010101001110110100: oled_data = 16'b1101111010011001;
				18'b010101010000110100: oled_data = 16'b1101111010111001;
				18'b010101010010110100: oled_data = 16'b1101011001111000;
				18'b010101010100110100: oled_data = 16'b1101011000010111;
				18'b010101010110110100: oled_data = 16'b1011110010010010;
				18'b010101011000110100: oled_data = 16'b1011001110101111;
				18'b010101011010110100: oled_data = 16'b1011101111010000;
				18'b010101011100110100: oled_data = 16'b1100010000110001;
				18'b010101011110110100: oled_data = 16'b1100110001010010;
				18'b010101100000110100: oled_data = 16'b1100010001010010;
				18'b010101100010110100: oled_data = 16'b1100010000010001;
				18'b010101100100110100: oled_data = 16'b1100110001110010;
				18'b010101100110110100: oled_data = 16'b1101010011010100;
				18'b010101101000110100: oled_data = 16'b1101010011010100;
				18'b010101101010110100: oled_data = 16'b1101010011010100;
				18'b010101101100110100: oled_data = 16'b1100110010010011;
				18'b010101101110110100: oled_data = 16'b1100010001110011;
				18'b010101110000110100: oled_data = 16'b1100010010010011;
				18'b010101110010110100: oled_data = 16'b1100010010010010;
				18'b010101110100110100: oled_data = 16'b1100010011010011;
				18'b010101110110110100: oled_data = 16'b1100110100110100;
				18'b010101111000110100: oled_data = 16'b1101010100010100;
				18'b010101111010110100: oled_data = 16'b1101010010110100;
				18'b010101111100110100: oled_data = 16'b1101010011010100;
				18'b010101111110110100: oled_data = 16'b1011001011101100;
				18'b010110000000110100: oled_data = 16'b1011001000001001;
				18'b010110000010110100: oled_data = 16'b1011001011001011;
				18'b010110000100110100: oled_data = 16'b1010101000001000;
				18'b010110000110110100: oled_data = 16'b1010101000001000;
				18'b010110001000110100: oled_data = 16'b1010101000001000;
				18'b010110001010110100: oled_data = 16'b1010101000001000;
				18'b010110001100110100: oled_data = 16'b1010101000001000;
				18'b010110001110110100: oled_data = 16'b1010101000001000;
				18'b010110010000110100: oled_data = 16'b1001101001001010;
				18'b010110010010110100: oled_data = 16'b1011111000011000;
				18'b010110010100110100: oled_data = 16'b1001111000111000;
				18'b010110010110110100: oled_data = 16'b1000110110010111;
				18'b010110011000110100: oled_data = 16'b1000110110010111;
				18'b010110011010110100: oled_data = 16'b1001010110110111;
				18'b010110011100110100: oled_data = 16'b1010001110101111;
				18'b010110011110110100: oled_data = 16'b1001100110100111;
				18'b010110100000110100: oled_data = 16'b1010000111000111;
				18'b010110100010110100: oled_data = 16'b1001100111000111;
				18'b010110100100110100: oled_data = 16'b1001100110100111;
				18'b010110100110110100: oled_data = 16'b1001100110100111;
				18'b010100011000110101: oled_data = 16'b1100001111110010;
				18'b010100011010110101: oled_data = 16'b1100001111110010;
				18'b010100011100110101: oled_data = 16'b1010001011001110;
				18'b010100011110110101: oled_data = 16'b1001101010001101;
				18'b010100100000110101: oled_data = 16'b1001101010101101;
				18'b010100100010110101: oled_data = 16'b1001101010101101;
				18'b010100100100110101: oled_data = 16'b1011001101110000;
				18'b010100100110110101: oled_data = 16'b1100110000010011;
				18'b010100101000110101: oled_data = 16'b1011001101110000;
				18'b010100101010110101: oled_data = 16'b1010001011001110;
				18'b010100101100110101: oled_data = 16'b1100001111110010;
				18'b010100101110110101: oled_data = 16'b1100010000010011;
				18'b010100110000110101: oled_data = 16'b1100110000010011;
				18'b010100110010110101: oled_data = 16'b1011101110110010;
				18'b010100110100110101: oled_data = 16'b1100001111010010;
				18'b010100110110110101: oled_data = 16'b1100110000010011;
				18'b010100111000110101: oled_data = 16'b1011001110010000;
				18'b010100111010110101: oled_data = 16'b1100010000010001;
				18'b010100111100110101: oled_data = 16'b1100010000010001;
				18'b010100111110110101: oled_data = 16'b1011101110110000;
				18'b010101000000110101: oled_data = 16'b1010101101101111;
				18'b010101000010110101: oled_data = 16'b1100110110010101;
				18'b010101000100110101: oled_data = 16'b1101111010011001;
				18'b010101000110110101: oled_data = 16'b1101111010011000;
				18'b010101001000110101: oled_data = 16'b1101111010011000;
				18'b010101001010110101: oled_data = 16'b1101111010011000;
				18'b010101001100110101: oled_data = 16'b1101111010011000;
				18'b010101001110110101: oled_data = 16'b1101111010011000;
				18'b010101010000110101: oled_data = 16'b1101111010011000;
				18'b010101010010110101: oled_data = 16'b1101111010011000;
				18'b010101010100110101: oled_data = 16'b1101011000110111;
				18'b010101010110110101: oled_data = 16'b1100110100110100;
				18'b010101011000110101: oled_data = 16'b1101010010110011;
				18'b010101011010110101: oled_data = 16'b1101010010110011;
				18'b010101011100110101: oled_data = 16'b1100110010110011;
				18'b010101011110110101: oled_data = 16'b1100110010010011;
				18'b010101100000110101: oled_data = 16'b1100110001110010;
				18'b010101100010110101: oled_data = 16'b1100010000110001;
				18'b010101100100110101: oled_data = 16'b1101010010110011;
				18'b010101100110110101: oled_data = 16'b1101010010110011;
				18'b010101101000110101: oled_data = 16'b1100110010010100;
				18'b010101101010110101: oled_data = 16'b1101010010010100;
				18'b010101101100110101: oled_data = 16'b1101010010010100;
				18'b010101101110110101: oled_data = 16'b1100010000110001;
				18'b010101110000110101: oled_data = 16'b1100010000110001;
				18'b010101110010110101: oled_data = 16'b1100110010010011;
				18'b010101110100110101: oled_data = 16'b1100110010010100;
				18'b010101110110110101: oled_data = 16'b1101010010010100;
				18'b010101111000110101: oled_data = 16'b1101010010010100;
				18'b010101111010110101: oled_data = 16'b1100110010010011;
				18'b010101111100110101: oled_data = 16'b1100010001010010;
				18'b010101111110110101: oled_data = 16'b1010001010001011;
				18'b010110000000110101: oled_data = 16'b1010100111101000;
				18'b010110000010110101: oled_data = 16'b1011001010001010;
				18'b010110000100110101: oled_data = 16'b1010101000001000;
				18'b010110000110110101: oled_data = 16'b1010101000001000;
				18'b010110001000110101: oled_data = 16'b1010101000001000;
				18'b010110001010110101: oled_data = 16'b1010101000001000;
				18'b010110001100110101: oled_data = 16'b1010100111101000;
				18'b010110001110110101: oled_data = 16'b1010000111101000;
				18'b010110010000110101: oled_data = 16'b1000100101000110;
				18'b010110010010110101: oled_data = 16'b1010101011001100;
				18'b010110010100110101: oled_data = 16'b1011010011010011;
				18'b010110010110110101: oled_data = 16'b1010010011010100;
				18'b010110011000110101: oled_data = 16'b1010010001010010;
				18'b010110011010110101: oled_data = 16'b1010001101001110;
				18'b010110011100110101: oled_data = 16'b1001100111101000;
				18'b010110011110110101: oled_data = 16'b1010000111000111;
				18'b010110100000110101: oled_data = 16'b1001100111000111;
				18'b010110100010110101: oled_data = 16'b1001100110100111;
				18'b010110100100110101: oled_data = 16'b1001100110100111;
				18'b010110100110110101: oled_data = 16'b1001100110100111;
				18'b010100011000110110: oled_data = 16'b1011101110110010;
				18'b010100011010110110: oled_data = 16'b1100001111010010;
				18'b010100011100110110: oled_data = 16'b1001101011001110;
				18'b010100011110110110: oled_data = 16'b1001001010001101;
				18'b010100100000110110: oled_data = 16'b1001101010001101;
				18'b010100100010110110: oled_data = 16'b1001001010001101;
				18'b010100100100110110: oled_data = 16'b1011001101010000;
				18'b010100100110110110: oled_data = 16'b1100001111110010;
				18'b010100101000110110: oled_data = 16'b1011001101010000;
				18'b010100101010110110: oled_data = 16'b1001101010001101;
				18'b010100101100110110: oled_data = 16'b1011101110010001;
				18'b010100101110110110: oled_data = 16'b1100001111110010;
				18'b010100110000110110: oled_data = 16'b1100001111010010;
				18'b010100110010110110: oled_data = 16'b1100001110110010;
				18'b010100110100110110: oled_data = 16'b1011101110110001;
				18'b010100110110110110: oled_data = 16'b1100110000010011;
				18'b010100111000110110: oled_data = 16'b1011001110010000;
				18'b010100111010110110: oled_data = 16'b1100010001010010;
				18'b010100111100110110: oled_data = 16'b1101010010110100;
				18'b010100111110110110: oled_data = 16'b1100110001010011;
				18'b010101000000110110: oled_data = 16'b1100010010010011;
				18'b010101000010110110: oled_data = 16'b1101011001011000;
				18'b010101000100110110: oled_data = 16'b1101011001111000;
				18'b010101000110110110: oled_data = 16'b1101011001111000;
				18'b010101001000110110: oled_data = 16'b1101011001111000;
				18'b010101001010110110: oled_data = 16'b1101011001111000;
				18'b010101001100110110: oled_data = 16'b1101011001111000;
				18'b010101001110110110: oled_data = 16'b1101011001011000;
				18'b010101010000110110: oled_data = 16'b1101011001011000;
				18'b010101010010110110: oled_data = 16'b1101011001011000;
				18'b010101010100110110: oled_data = 16'b1101011001011000;
				18'b010101010110110110: oled_data = 16'b1100110100110101;
				18'b010101011000110110: oled_data = 16'b1100110001110011;
				18'b010101011010110110: oled_data = 16'b1100110010010011;
				18'b010101011100110110: oled_data = 16'b1100110010010011;
				18'b010101011110110110: oled_data = 16'b1100110010010011;
				18'b010101100000110110: oled_data = 16'b1100110010010011;
				18'b010101100010110110: oled_data = 16'b1100010000110001;
				18'b010101100100110110: oled_data = 16'b1100110001110010;
				18'b010101100110110110: oled_data = 16'b1100110001110011;
				18'b010101101000110110: oled_data = 16'b1100110001110011;
				18'b010101101010110110: oled_data = 16'b1100110001110011;
				18'b010101101100110110: oled_data = 16'b1100110001110011;
				18'b010101101110110110: oled_data = 16'b1100110001110010;
				18'b010101110000110110: oled_data = 16'b1100010000110001;
				18'b010101110010110110: oled_data = 16'b1011001111010001;
				18'b010101110100110110: oled_data = 16'b1100010000110010;
				18'b010101110110110110: oled_data = 16'b1100110001010011;
				18'b010101111000110110: oled_data = 16'b1100010000110010;
				18'b010101111010110110: oled_data = 16'b1100010000110001;
				18'b010101111100110110: oled_data = 16'b1100010001010010;
				18'b010101111110110110: oled_data = 16'b1010001010101011;
				18'b010110000000110110: oled_data = 16'b1010100111101000;
				18'b010110000010110110: oled_data = 16'b1010101001101001;
				18'b010110000100110110: oled_data = 16'b1010100111101000;
				18'b010110000110110110: oled_data = 16'b1010100111101000;
				18'b010110001000110110: oled_data = 16'b1010100111101000;
				18'b010110001010110110: oled_data = 16'b1010000111101000;
				18'b010110001100110110: oled_data = 16'b1010100111100111;
				18'b010110001110110110: oled_data = 16'b1001100111000111;
				18'b010110010000110110: oled_data = 16'b1000100110000110;
				18'b010110010010110110: oled_data = 16'b1010000111000111;
				18'b010110010100110110: oled_data = 16'b1010000111000111;
				18'b010110010110110110: oled_data = 16'b1010000111101000;
				18'b010110011000110110: oled_data = 16'b1001100110100111;
				18'b010110011010110110: oled_data = 16'b1010000110100111;
				18'b010110011100110110: oled_data = 16'b1001100111000111;
				18'b010110011110110110: oled_data = 16'b1001100110100111;
				18'b010110100000110110: oled_data = 16'b1001100110100111;
				18'b010110100010110110: oled_data = 16'b1001100110100110;
				18'b010110100100110110: oled_data = 16'b1001000110000110;
				18'b010110100110110110: oled_data = 16'b1001000110000110;
				18'b010100011000110111: oled_data = 16'b1100001110110001;
				18'b010100011010110111: oled_data = 16'b1100001110110001;
				18'b010100011100110111: oled_data = 16'b1001101010101101;
				18'b010100011110110111: oled_data = 16'b1001001010001101;
				18'b010100100000110111: oled_data = 16'b1001001010001101;
				18'b010100100010110111: oled_data = 16'b1001001010001101;
				18'b010100100100110111: oled_data = 16'b1011001101010000;
				18'b010100100110110111: oled_data = 16'b1100001111010010;
				18'b010100101000110111: oled_data = 16'b1011001101110000;
				18'b010100101010110111: oled_data = 16'b1001001010001101;
				18'b010100101100110111: oled_data = 16'b1011001101010000;
				18'b010100101110110111: oled_data = 16'b1100001110110001;
				18'b010100110000110111: oled_data = 16'b1100001110110010;
				18'b010100110010110111: oled_data = 16'b1011101110010001;
				18'b010100110100110111: oled_data = 16'b1011101110010001;
				18'b010100110110110111: oled_data = 16'b1100001111010010;
				18'b010100111000110111: oled_data = 16'b1011101110110001;
				18'b010100111010110111: oled_data = 16'b1100001111110010;
				18'b010100111100110111: oled_data = 16'b1100110001010011;
				18'b010100111110110111: oled_data = 16'b1100001111110010;
				18'b010101000000110111: oled_data = 16'b1100110011110100;
				18'b010101000010110111: oled_data = 16'b1101011001011000;
				18'b010101000100110111: oled_data = 16'b1101011001010111;
				18'b010101000110110111: oled_data = 16'b1101011001010111;
				18'b010101001000110111: oled_data = 16'b1101011001010111;
				18'b010101001010110111: oled_data = 16'b1101011000110111;
				18'b010101001100110111: oled_data = 16'b1101011000110111;
				18'b010101001110110111: oled_data = 16'b1101011000110111;
				18'b010101010000110111: oled_data = 16'b1101011000110111;
				18'b010101010010110111: oled_data = 16'b1101011000110111;
				18'b010101010100110111: oled_data = 16'b1101011000010111;
				18'b010101010110110111: oled_data = 16'b1100010010110011;
				18'b010101011000110111: oled_data = 16'b1100110001010010;
				18'b010101011010110111: oled_data = 16'b1100110001010010;
				18'b010101011100110111: oled_data = 16'b1100110001110010;
				18'b010101011110110111: oled_data = 16'b1100110001110010;
				18'b010101100000110111: oled_data = 16'b1100110001110010;
				18'b010101100010110111: oled_data = 16'b1100010000010001;
				18'b010101100100110111: oled_data = 16'b1100110001010010;
				18'b010101100110110111: oled_data = 16'b1100110001010010;
				18'b010101101000110111: oled_data = 16'b1100110001010010;
				18'b010101101010110111: oled_data = 16'b1100110001010010;
				18'b010101101100110111: oled_data = 16'b1100110001010010;
				18'b010101101110110111: oled_data = 16'b1100110001110011;
				18'b010101110000110111: oled_data = 16'b1011110000010001;
				18'b010101110010110111: oled_data = 16'b0110000110100111;
				18'b010101110100110111: oled_data = 16'b1011001111010000;
				18'b010101110110110111: oled_data = 16'b1100010000110010;
				18'b010101111000110111: oled_data = 16'b1100010000110001;
				18'b010101111010110111: oled_data = 16'b1100110001110010;
				18'b010101111100110111: oled_data = 16'b1100110001110011;
				18'b010101111110110111: oled_data = 16'b1010001010101100;
				18'b010110000000110111: oled_data = 16'b1010100111100111;
				18'b010110000010110111: oled_data = 16'b1010001000101000;
				18'b010110000100110111: oled_data = 16'b1010100111101000;
				18'b010110000110110111: oled_data = 16'b1010100111100111;
				18'b010110001000110111: oled_data = 16'b1010000111100111;
				18'b010110001010110111: oled_data = 16'b1010000111100111;
				18'b010110001100110111: oled_data = 16'b1010000111000111;
				18'b010110001110110111: oled_data = 16'b1001100110100111;
				18'b010110010000110111: oled_data = 16'b1000100110000111;
				18'b010110010010110111: oled_data = 16'b1010000111001000;
				18'b010110010100110111: oled_data = 16'b1010000111000111;
				18'b010110010110110111: oled_data = 16'b1001100110100111;
				18'b010110011000110111: oled_data = 16'b1001000110100110;
				18'b010110011010110111: oled_data = 16'b1001100110100111;
				18'b010110011100110111: oled_data = 16'b1001100110100111;
				18'b010110011110110111: oled_data = 16'b1001100110100110;
				18'b010110100000110111: oled_data = 16'b1001100110000110;
				18'b010110100010110111: oled_data = 16'b1001000110000110;
				18'b010110100100110111: oled_data = 16'b1001000110000110;
				18'b010110100110110111: oled_data = 16'b1001000110000110;
				18'b011000011000001000: oled_data = 16'b1001101111101011;
				18'b011000011010001000: oled_data = 16'b1010010000001011;
				18'b011000011100001000: oled_data = 16'b1010010000101011;
				18'b011000011110001000: oled_data = 16'b1010110000101011;
				18'b011000100000001000: oled_data = 16'b1011010001101101;
				18'b011000100010001000: oled_data = 16'b1110011000111000;
				18'b011000100100001000: oled_data = 16'b1110010101010111;
				18'b011000100110001000: oled_data = 16'b1101110011010101;
				18'b011000101000001000: oled_data = 16'b1101110011010101;
				18'b011000101010001000: oled_data = 16'b1101110011010101;
				18'b011000101100001000: oled_data = 16'b1101110011010101;
				18'b011000101110001000: oled_data = 16'b1101110011010101;
				18'b011000110000001000: oled_data = 16'b1101110011010101;
				18'b011000110010001000: oled_data = 16'b1101110011010101;
				18'b011000110100001000: oled_data = 16'b1101110011010101;
				18'b011000110110001000: oled_data = 16'b1101110011010101;
				18'b011000111000001000: oled_data = 16'b1101110011010101;
				18'b011000111010001000: oled_data = 16'b1101110011010101;
				18'b011000111100001000: oled_data = 16'b1101110011010101;
				18'b011000111110001000: oled_data = 16'b1101110011010101;
				18'b011001000000001000: oled_data = 16'b1101110011010101;
				18'b011001000010001000: oled_data = 16'b1101110011010101;
				18'b011001000100001000: oled_data = 16'b1101110011010101;
				18'b011001000110001000: oled_data = 16'b1101110011010101;
				18'b011001001000001000: oled_data = 16'b1101110011010101;
				18'b011001001010001000: oled_data = 16'b1101110011010101;
				18'b011001001100001000: oled_data = 16'b1101110011010101;
				18'b011001001110001000: oled_data = 16'b1101110011010101;
				18'b011001010000001000: oled_data = 16'b1101110011010101;
				18'b011001010010001000: oled_data = 16'b1101110011010101;
				18'b011001010100001000: oled_data = 16'b1101110011010101;
				18'b011001010110001000: oled_data = 16'b1101110011010101;
				18'b011001011000001000: oled_data = 16'b1101110011010101;
				18'b011001011010001000: oled_data = 16'b1101110011010101;
				18'b011001011100001000: oled_data = 16'b1101110011010101;
				18'b011001011110001000: oled_data = 16'b1101110011010101;
				18'b011001100000001000: oled_data = 16'b1101110011010101;
				18'b011001100010001000: oled_data = 16'b1101110011010101;
				18'b011001100100001000: oled_data = 16'b1101110011010101;
				18'b011001100110001000: oled_data = 16'b1101110011010101;
				18'b011001101000001000: oled_data = 16'b1101110011010101;
				18'b011001101010001000: oled_data = 16'b1101110011010101;
				18'b011001101100001000: oled_data = 16'b1101110011010101;
				18'b011001101110001000: oled_data = 16'b1101110011010101;
				18'b011001110000001000: oled_data = 16'b1101110011010101;
				18'b011001110010001000: oled_data = 16'b1101110100010110;
				18'b011001110100001000: oled_data = 16'b1110111000111010;
				18'b011001110110001000: oled_data = 16'b1011110110010110;
				18'b011001111000001000: oled_data = 16'b1010010100110100;
				18'b011001111010001000: oled_data = 16'b1010010101010100;
				18'b011001111100001000: oled_data = 16'b0101101011001011;
				18'b011001111110001000: oled_data = 16'b0100001000001000;
				18'b011010000000001000: oled_data = 16'b0100001000101000;
				18'b011010000010001000: oled_data = 16'b0100001000101000;
				18'b011010000100001000: oled_data = 16'b0100001000100111;
				18'b011010000110001000: oled_data = 16'b0011100110100110;
				18'b011010001000001000: oled_data = 16'b0101000111100101;
				18'b011010001010001000: oled_data = 16'b0110001001000101;
				18'b011010001100001000: oled_data = 16'b0111001011000111;
				18'b011010001110001000: oled_data = 16'b0111101100001000;
				18'b011010010000001000: oled_data = 16'b0111101100001000;
				18'b011010010010001000: oled_data = 16'b0111101100001000;
				18'b011010010100001000: oled_data = 16'b0111101100001000;
				18'b011010010110001000: oled_data = 16'b0111001011101000;
				18'b011010011000001000: oled_data = 16'b0110101011101000;
				18'b011010011010001000: oled_data = 16'b0110001011001000;
				18'b011010011100001000: oled_data = 16'b0110001010101000;
				18'b011010011110001000: oled_data = 16'b0101101010001000;
				18'b011010100000001000: oled_data = 16'b0101101010001000;
				18'b011010100010001000: oled_data = 16'b0101001001101000;
				18'b011010100100001000: oled_data = 16'b0101001001001000;
				18'b011010100110001000: oled_data = 16'b0101001001101000;
				18'b011000011000001001: oled_data = 16'b1011010001101100;
				18'b011000011010001001: oled_data = 16'b1011010001001011;
				18'b011000011100001001: oled_data = 16'b1011010001001011;
				18'b011000011110001001: oled_data = 16'b1010110000101011;
				18'b011000100000001001: oled_data = 16'b1101010110010100;
				18'b011000100010001001: oled_data = 16'b1110010110011000;
				18'b011000100100001001: oled_data = 16'b1101110011010110;
				18'b011000100110001001: oled_data = 16'b1101110011010101;
				18'b011000101000001001: oled_data = 16'b1101110011010101;
				18'b011000101010001001: oled_data = 16'b1101110011010101;
				18'b011000101100001001: oled_data = 16'b1101110011010101;
				18'b011000101110001001: oled_data = 16'b1101110011010101;
				18'b011000110000001001: oled_data = 16'b1101110011010101;
				18'b011000110010001001: oled_data = 16'b1101110011010101;
				18'b011000110100001001: oled_data = 16'b1101110011010101;
				18'b011000110110001001: oled_data = 16'b1101110011010101;
				18'b011000111000001001: oled_data = 16'b1101110011010101;
				18'b011000111010001001: oled_data = 16'b1101110011010101;
				18'b011000111100001001: oled_data = 16'b1101110011010101;
				18'b011000111110001001: oled_data = 16'b1101110011010101;
				18'b011001000000001001: oled_data = 16'b1101110011010101;
				18'b011001000010001001: oled_data = 16'b1101110011010101;
				18'b011001000100001001: oled_data = 16'b1101110011010101;
				18'b011001000110001001: oled_data = 16'b1101110011010101;
				18'b011001001000001001: oled_data = 16'b1101110011010101;
				18'b011001001010001001: oled_data = 16'b1101110011010101;
				18'b011001001100001001: oled_data = 16'b1101110011010101;
				18'b011001001110001001: oled_data = 16'b1101110011010101;
				18'b011001010000001001: oled_data = 16'b1101110011010101;
				18'b011001010010001001: oled_data = 16'b1101110011010101;
				18'b011001010100001001: oled_data = 16'b1101110011010101;
				18'b011001010110001001: oled_data = 16'b1101110011010101;
				18'b011001011000001001: oled_data = 16'b1101110011010101;
				18'b011001011010001001: oled_data = 16'b1101110011010101;
				18'b011001011100001001: oled_data = 16'b1101110011010101;
				18'b011001011110001001: oled_data = 16'b1101110011010101;
				18'b011001100000001001: oled_data = 16'b1101110011010101;
				18'b011001100010001001: oled_data = 16'b1101110011010101;
				18'b011001100100001001: oled_data = 16'b1101110011010101;
				18'b011001100110001001: oled_data = 16'b1101110011010101;
				18'b011001101000001001: oled_data = 16'b1101110011010101;
				18'b011001101010001001: oled_data = 16'b1101110011010101;
				18'b011001101100001001: oled_data = 16'b1101110011010101;
				18'b011001101110001001: oled_data = 16'b1101110011010101;
				18'b011001110000001001: oled_data = 16'b1101110011010101;
				18'b011001110010001001: oled_data = 16'b1101110010110101;
				18'b011001110100001001: oled_data = 16'b1110010101010111;
				18'b011001110110001001: oled_data = 16'b1110111001111010;
				18'b011001111000001001: oled_data = 16'b1010010011010011;
				18'b011001111010001001: oled_data = 16'b0111001110001110;
				18'b011001111100001001: oled_data = 16'b0100101001101001;
				18'b011001111110001001: oled_data = 16'b0100001000001000;
				18'b011010000000001001: oled_data = 16'b0100001000101000;
				18'b011010000010001001: oled_data = 16'b0100001000101000;
				18'b011010000100001001: oled_data = 16'b0100001000000111;
				18'b011010000110001001: oled_data = 16'b0011100110100101;
				18'b011010001000001001: oled_data = 16'b0100100110100100;
				18'b011010001010001001: oled_data = 16'b0101101000100101;
				18'b011010001100001001: oled_data = 16'b0111001010100111;
				18'b011010001110001001: oled_data = 16'b0111101100001000;
				18'b011010010000001001: oled_data = 16'b1000001100101000;
				18'b011010010010001001: oled_data = 16'b1000001100101000;
				18'b011010010100001001: oled_data = 16'b1000001100101000;
				18'b011010010110001001: oled_data = 16'b1000001101001000;
				18'b011010011000001001: oled_data = 16'b1000101101101000;
				18'b011010011010001001: oled_data = 16'b1000101101101000;
				18'b011010011100001001: oled_data = 16'b1000101101101000;
				18'b011010011110001001: oled_data = 16'b1000101110001001;
				18'b011010100000001001: oled_data = 16'b1000101110101001;
				18'b011010100010001001: oled_data = 16'b0101101010101000;
				18'b011010100100001001: oled_data = 16'b0011101000000111;
				18'b011010100110001001: oled_data = 16'b0100001000001000;
				18'b011000011000001010: oled_data = 16'b1011010001101100;
				18'b011000011010001010: oled_data = 16'b1011010001101011;
				18'b011000011100001010: oled_data = 16'b1010110001001011;
				18'b011000011110001010: oled_data = 16'b1100010010110000;
				18'b011000100000001010: oled_data = 16'b1110010101010110;
				18'b011000100010001010: oled_data = 16'b1101110010110101;
				18'b011000100100001010: oled_data = 16'b1101110011010110;
				18'b011000100110001010: oled_data = 16'b1101110011010101;
				18'b011000101000001010: oled_data = 16'b1101110011010101;
				18'b011000101010001010: oled_data = 16'b1101110011010101;
				18'b011000101100001010: oled_data = 16'b1101110011010101;
				18'b011000101110001010: oled_data = 16'b1101110011010101;
				18'b011000110000001010: oled_data = 16'b1101110011010101;
				18'b011000110010001010: oled_data = 16'b1101110011010101;
				18'b011000110100001010: oled_data = 16'b1101110011010101;
				18'b011000110110001010: oled_data = 16'b1101110011010101;
				18'b011000111000001010: oled_data = 16'b1101110011010101;
				18'b011000111010001010: oled_data = 16'b1101110011010101;
				18'b011000111100001010: oled_data = 16'b1101110011010101;
				18'b011000111110001010: oled_data = 16'b1101110011010101;
				18'b011001000000001010: oled_data = 16'b1101110011010101;
				18'b011001000010001010: oled_data = 16'b1101110011010101;
				18'b011001000100001010: oled_data = 16'b1101110011010101;
				18'b011001000110001010: oled_data = 16'b1101110011010101;
				18'b011001001000001010: oled_data = 16'b1101110011010101;
				18'b011001001010001010: oled_data = 16'b1101110011010101;
				18'b011001001100001010: oled_data = 16'b1101110011010101;
				18'b011001001110001010: oled_data = 16'b1101110011010101;
				18'b011001010000001010: oled_data = 16'b1101110011010101;
				18'b011001010010001010: oled_data = 16'b1101110011010101;
				18'b011001010100001010: oled_data = 16'b1101110011010101;
				18'b011001010110001010: oled_data = 16'b1101110011010101;
				18'b011001011000001010: oled_data = 16'b1101110011010101;
				18'b011001011010001010: oled_data = 16'b1101110011010101;
				18'b011001011100001010: oled_data = 16'b1101110011010101;
				18'b011001011110001010: oled_data = 16'b1101110011010101;
				18'b011001100000001010: oled_data = 16'b1101110011010101;
				18'b011001100010001010: oled_data = 16'b1101110011010101;
				18'b011001100100001010: oled_data = 16'b1101110011010101;
				18'b011001100110001010: oled_data = 16'b1101110011010101;
				18'b011001101000001010: oled_data = 16'b1101110011010110;
				18'b011001101010001010: oled_data = 16'b1110010011010110;
				18'b011001101100001010: oled_data = 16'b1110010011010110;
				18'b011001101110001010: oled_data = 16'b1110010011010110;
				18'b011001110000001010: oled_data = 16'b1110010011010110;
				18'b011001110010001010: oled_data = 16'b1101110011010101;
				18'b011001110100001010: oled_data = 16'b1101110011010101;
				18'b011001110110001010: oled_data = 16'b1110110110011000;
				18'b011001111000001010: oled_data = 16'b1100110101010110;
				18'b011001111010001010: oled_data = 16'b0101001000101001;
				18'b011001111100001010: oled_data = 16'b0100001000001000;
				18'b011001111110001010: oled_data = 16'b0011101000000111;
				18'b011010000000001010: oled_data = 16'b0011100111100111;
				18'b011010000010001010: oled_data = 16'b0100001000101000;
				18'b011010000100001010: oled_data = 16'b0100001000101000;
				18'b011010000110001010: oled_data = 16'b0011000101100101;
				18'b011010001000001010: oled_data = 16'b0010100100100100;
				18'b011010001010001010: oled_data = 16'b0011000101100101;
				18'b011010001100001010: oled_data = 16'b0100000111000110;
				18'b011010001110001010: oled_data = 16'b0101001000100110;
				18'b011010010000001010: oled_data = 16'b0110001010000111;
				18'b011010010010001010: oled_data = 16'b0111001011001000;
				18'b011010010100001010: oled_data = 16'b0111001011101000;
				18'b011010010110001010: oled_data = 16'b0111101100001000;
				18'b011010011000001010: oled_data = 16'b1000101101001000;
				18'b011010011010001010: oled_data = 16'b1000101101101000;
				18'b011010011100001010: oled_data = 16'b1000101110001000;
				18'b011010011110001010: oled_data = 16'b1001001110001000;
				18'b011010100000001010: oled_data = 16'b1000101110001001;
				18'b011010100010001010: oled_data = 16'b0111001011101001;
				18'b011010100100001010: oled_data = 16'b1001001101001101;
				18'b011010100110001010: oled_data = 16'b1011010000110001;
				18'b011000011000001011: oled_data = 16'b1001001111001010;
				18'b011000011010001011: oled_data = 16'b1000101101101001;
				18'b011000011100001011: oled_data = 16'b1001001111001100;
				18'b011000011110001011: oled_data = 16'b1101010100110101;
				18'b011000100000001011: oled_data = 16'b1101010010010100;
				18'b011000100010001011: oled_data = 16'b1101110010110101;
				18'b011000100100001011: oled_data = 16'b1101110011010101;
				18'b011000100110001011: oled_data = 16'b1101110010110101;
				18'b011000101000001011: oled_data = 16'b1101010010010100;
				18'b011000101010001011: oled_data = 16'b1101110011010110;
				18'b011000101100001011: oled_data = 16'b1101110011010101;
				18'b011000101110001011: oled_data = 16'b1101110011010101;
				18'b011000110000001011: oled_data = 16'b1101110011010101;
				18'b011000110010001011: oled_data = 16'b1101110011010101;
				18'b011000110100001011: oled_data = 16'b1101110011010101;
				18'b011000110110001011: oled_data = 16'b1101110011010101;
				18'b011000111000001011: oled_data = 16'b1101110011010101;
				18'b011000111010001011: oled_data = 16'b1101110011010101;
				18'b011000111100001011: oled_data = 16'b1101110011010101;
				18'b011000111110001011: oled_data = 16'b1101110011010101;
				18'b011001000000001011: oled_data = 16'b1101110011010101;
				18'b011001000010001011: oled_data = 16'b1101110011010101;
				18'b011001000100001011: oled_data = 16'b1101110011010101;
				18'b011001000110001011: oled_data = 16'b1101110011010101;
				18'b011001001000001011: oled_data = 16'b1101110011010101;
				18'b011001001010001011: oled_data = 16'b1101110011010101;
				18'b011001001100001011: oled_data = 16'b1101110011010101;
				18'b011001001110001011: oled_data = 16'b1101110011010101;
				18'b011001010000001011: oled_data = 16'b1101110011010101;
				18'b011001010010001011: oled_data = 16'b1101110011010101;
				18'b011001010100001011: oled_data = 16'b1101110011010101;
				18'b011001010110001011: oled_data = 16'b1101110011010101;
				18'b011001011000001011: oled_data = 16'b1101110011010101;
				18'b011001011010001011: oled_data = 16'b1101110011010101;
				18'b011001011100001011: oled_data = 16'b1101110011010101;
				18'b011001011110001011: oled_data = 16'b1101110011010101;
				18'b011001100000001011: oled_data = 16'b1101110011010101;
				18'b011001100010001011: oled_data = 16'b1101110011010101;
				18'b011001100100001011: oled_data = 16'b1101110011010101;
				18'b011001100110001011: oled_data = 16'b1110010011010110;
				18'b011001101000001011: oled_data = 16'b1110010011010110;
				18'b011001101010001011: oled_data = 16'b1110010011010110;
				18'b011001101100001011: oled_data = 16'b1110010011010110;
				18'b011001101110001011: oled_data = 16'b1101110011010110;
				18'b011001110000001011: oled_data = 16'b1101110011010110;
				18'b011001110010001011: oled_data = 16'b1101110011010101;
				18'b011001110100001011: oled_data = 16'b1101110011010101;
				18'b011001110110001011: oled_data = 16'b1101110011110110;
				18'b011001111000001011: oled_data = 16'b1111010111111001;
				18'b011001111010001011: oled_data = 16'b1001001111110000;
				18'b011001111100001011: oled_data = 16'b0100001000000111;
				18'b011001111110001011: oled_data = 16'b0100101010001000;
				18'b011010000000001011: oled_data = 16'b0101101011001001;
				18'b011010000010001011: oled_data = 16'b0110001100101011;
				18'b011010000100001011: oled_data = 16'b0110001100001011;
				18'b011010000110001011: oled_data = 16'b0010100101100101;
				18'b011010001000001011: oled_data = 16'b0001100011100011;
				18'b011010001010001011: oled_data = 16'b0010000100100100;
				18'b011010001100001011: oled_data = 16'b0010000101000110;
				18'b011010001110001011: oled_data = 16'b0010000101000101;
				18'b011010010000001011: oled_data = 16'b0010100101100110;
				18'b011010010010001011: oled_data = 16'b0011000110000110;
				18'b011010010100001011: oled_data = 16'b0011100111000111;
				18'b011010010110001011: oled_data = 16'b0100000111100111;
				18'b011010011000001011: oled_data = 16'b0101001000100111;
				18'b011010011010001011: oled_data = 16'b0101101001100111;
				18'b011010011100001011: oled_data = 16'b0111001011001000;
				18'b011010011110001011: oled_data = 16'b1010001110001100;
				18'b011010100000001011: oled_data = 16'b1100010001010000;
				18'b011010100010001011: oled_data = 16'b1101110010110010;
				18'b011010100100001011: oled_data = 16'b1101110001010001;
				18'b011010100110001011: oled_data = 16'b1100101110001110;
				18'b011000011000001100: oled_data = 16'b0110001010001000;
				18'b011000011010001100: oled_data = 16'b0110001010001000;
				18'b011000011100001100: oled_data = 16'b1010110001010001;
				18'b011000011110001100: oled_data = 16'b1101010011010101;
				18'b011000100000001100: oled_data = 16'b1101110010010101;
				18'b011000100010001100: oled_data = 16'b1101110011010101;
				18'b011000100100001100: oled_data = 16'b1101110011010110;
				18'b011000100110001100: oled_data = 16'b1101010010010100;
				18'b011000101000001100: oled_data = 16'b1101110010110101;
				18'b011000101010001100: oled_data = 16'b1101110011010101;
				18'b011000101100001100: oled_data = 16'b1101110011010101;
				18'b011000101110001100: oled_data = 16'b1101110011010101;
				18'b011000110000001100: oled_data = 16'b1101110011010101;
				18'b011000110010001100: oled_data = 16'b1101110011010101;
				18'b011000110100001100: oled_data = 16'b1101110011010101;
				18'b011000110110001100: oled_data = 16'b1101110011010101;
				18'b011000111000001100: oled_data = 16'b1101110011010101;
				18'b011000111010001100: oled_data = 16'b1101110011010101;
				18'b011000111100001100: oled_data = 16'b1101110011010101;
				18'b011000111110001100: oled_data = 16'b1101110011010101;
				18'b011001000000001100: oled_data = 16'b1101110010110101;
				18'b011001000010001100: oled_data = 16'b1101110011010101;
				18'b011001000100001100: oled_data = 16'b1101110011010101;
				18'b011001000110001100: oled_data = 16'b1101110011010101;
				18'b011001001000001100: oled_data = 16'b1101110011010101;
				18'b011001001010001100: oled_data = 16'b1101110011010101;
				18'b011001001100001100: oled_data = 16'b1101110011010101;
				18'b011001001110001100: oled_data = 16'b1101110011010101;
				18'b011001010000001100: oled_data = 16'b1101110011010101;
				18'b011001010010001100: oled_data = 16'b1101110011010101;
				18'b011001010100001100: oled_data = 16'b1101110011010101;
				18'b011001010110001100: oled_data = 16'b1101110011010101;
				18'b011001011000001100: oled_data = 16'b1101110011010101;
				18'b011001011010001100: oled_data = 16'b1101110011010101;
				18'b011001011100001100: oled_data = 16'b1101110011010101;
				18'b011001011110001100: oled_data = 16'b1101110011010101;
				18'b011001100000001100: oled_data = 16'b1101110011010101;
				18'b011001100010001100: oled_data = 16'b1101110011010101;
				18'b011001100100001100: oled_data = 16'b1101110011010101;
				18'b011001100110001100: oled_data = 16'b1101110011010110;
				18'b011001101000001100: oled_data = 16'b1110010011010110;
				18'b011001101010001100: oled_data = 16'b1101110011010110;
				18'b011001101100001100: oled_data = 16'b1101110011010110;
				18'b011001101110001100: oled_data = 16'b1101110011010101;
				18'b011001110000001100: oled_data = 16'b1101110011010101;
				18'b011001110010001100: oled_data = 16'b1101110011010110;
				18'b011001110100001100: oled_data = 16'b1101110011010110;
				18'b011001110110001100: oled_data = 16'b1101110011010101;
				18'b011001111000001100: oled_data = 16'b1110010100010110;
				18'b011001111010001100: oled_data = 16'b1101110110111000;
				18'b011001111100001100: oled_data = 16'b0111001101001011;
				18'b011001111110001100: oled_data = 16'b0110101101001001;
				18'b011010000000001100: oled_data = 16'b0111101110101011;
				18'b011010000010001100: oled_data = 16'b1000010000001100;
				18'b011010000100001100: oled_data = 16'b0110101101101011;
				18'b011010000110001100: oled_data = 16'b0010000100100100;
				18'b011010001000001100: oled_data = 16'b0001100011000011;
				18'b011010001010001100: oled_data = 16'b0001100100000100;
				18'b011010001100001100: oled_data = 16'b0010000100100101;
				18'b011010001110001100: oled_data = 16'b0010000101000101;
				18'b011010010000001100: oled_data = 16'b0010000101000110;
				18'b011010010010001100: oled_data = 16'b0010100101100110;
				18'b011010010100001100: oled_data = 16'b0010100110000111;
				18'b011010010110001100: oled_data = 16'b0010100110000111;
				18'b011010011000001100: oled_data = 16'b0010100110100111;
				18'b011010011010001100: oled_data = 16'b0110101010101011;
				18'b011010011100001100: oled_data = 16'b1011110001010001;
				18'b011010011110001100: oled_data = 16'b1110010011010011;
				18'b011010100000001100: oled_data = 16'b1101110000110001;
				18'b011010100010001100: oled_data = 16'b1100001100001100;
				18'b011010100100001100: oled_data = 16'b1010101001001001;
				18'b011010100110001100: oled_data = 16'b1010101000001000;
				18'b011000011000001101: oled_data = 16'b1000110001110000;
				18'b011000011010001101: oled_data = 16'b1001010010010000;
				18'b011000011100001101: oled_data = 16'b1100010100010100;
				18'b011000011110001101: oled_data = 16'b1101010010010100;
				18'b011000100000001101: oled_data = 16'b1101110011010101;
				18'b011000100010001101: oled_data = 16'b1101110011010101;
				18'b011000100100001101: oled_data = 16'b1101110011010101;
				18'b011000100110001101: oled_data = 16'b1101010010010100;
				18'b011000101000001101: oled_data = 16'b1101110011010101;
				18'b011000101010001101: oled_data = 16'b1101110011010101;
				18'b011000101100001101: oled_data = 16'b1101110011010101;
				18'b011000101110001101: oled_data = 16'b1101110011010101;
				18'b011000110000001101: oled_data = 16'b1101110010110101;
				18'b011000110010001101: oled_data = 16'b1101110011010101;
				18'b011000110100001101: oled_data = 16'b1101110011010101;
				18'b011000110110001101: oled_data = 16'b1101110011010101;
				18'b011000111000001101: oled_data = 16'b1101110011010101;
				18'b011000111010001101: oled_data = 16'b1101110011010101;
				18'b011000111100001101: oled_data = 16'b1101110011010101;
				18'b011000111110001101: oled_data = 16'b1101110011010110;
				18'b011001000000001101: oled_data = 16'b1101110010010101;
				18'b011001000010001101: oled_data = 16'b1101110010110101;
				18'b011001000100001101: oled_data = 16'b1101110011010110;
				18'b011001000110001101: oled_data = 16'b1101110011010101;
				18'b011001001000001101: oled_data = 16'b1101110011010101;
				18'b011001001010001101: oled_data = 16'b1101110011010101;
				18'b011001001100001101: oled_data = 16'b1101110011010101;
				18'b011001001110001101: oled_data = 16'b1101110011010101;
				18'b011001010000001101: oled_data = 16'b1101110011010101;
				18'b011001010010001101: oled_data = 16'b1101110011010101;
				18'b011001010100001101: oled_data = 16'b1101110011010101;
				18'b011001010110001101: oled_data = 16'b1101110011010101;
				18'b011001011000001101: oled_data = 16'b1101110011010101;
				18'b011001011010001101: oled_data = 16'b1101110011010101;
				18'b011001011100001101: oled_data = 16'b1101110011010101;
				18'b011001011110001101: oled_data = 16'b1101110011010101;
				18'b011001100000001101: oled_data = 16'b1101110011010101;
				18'b011001100010001101: oled_data = 16'b1101110011010101;
				18'b011001100100001101: oled_data = 16'b1101110011010101;
				18'b011001100110001101: oled_data = 16'b1101110011010101;
				18'b011001101000001101: oled_data = 16'b1101110011010101;
				18'b011001101010001101: oled_data = 16'b1101110011010101;
				18'b011001101100001101: oled_data = 16'b1101110011010101;
				18'b011001101110001101: oled_data = 16'b1101110011010101;
				18'b011001110000001101: oled_data = 16'b1101110011010101;
				18'b011001110010001101: oled_data = 16'b1110010011010110;
				18'b011001110100001101: oled_data = 16'b1110010011010110;
				18'b011001110110001101: oled_data = 16'b1110010011010110;
				18'b011001111000001101: oled_data = 16'b1101110011010101;
				18'b011001111010001101: oled_data = 16'b1111010111011001;
				18'b011001111100001101: oled_data = 16'b1010110011010010;
				18'b011001111110001101: oled_data = 16'b0110001011101000;
				18'b011010000000001101: oled_data = 16'b0110101101001001;
				18'b011010000010001101: oled_data = 16'b0110101100101000;
				18'b011010000100001101: oled_data = 16'b0100101001100111;
				18'b011010000110001101: oled_data = 16'b0001100011000011;
				18'b011010001000001101: oled_data = 16'b0001100011000011;
				18'b011010001010001101: oled_data = 16'b0001100100000100;
				18'b011010001100001101: oled_data = 16'b0010000100100100;
				18'b011010001110001101: oled_data = 16'b0010000101000101;
				18'b011010010000001101: oled_data = 16'b0010000101000110;
				18'b011010010010001101: oled_data = 16'b0010000101000110;
				18'b011010010100001101: oled_data = 16'b0010000101000110;
				18'b011010010110001101: oled_data = 16'b0100001000001000;
				18'b011010011000001101: oled_data = 16'b1010101111110000;
				18'b011010011010001101: oled_data = 16'b1110010100010100;
				18'b011010011100001101: oled_data = 16'b1110010010010010;
				18'b011010011110001101: oled_data = 16'b1100001100101101;
				18'b011010100000001101: oled_data = 16'b1011001001001001;
				18'b011010100010001101: oled_data = 16'b1011001000001000;
				18'b011010100100001101: oled_data = 16'b1010101000101000;
				18'b011010100110001101: oled_data = 16'b1010101000001000;
				18'b011000011000001110: oled_data = 16'b0111111000111010;
				18'b011000011010001110: oled_data = 16'b1000110110110111;
				18'b011000011100001110: oled_data = 16'b1100110010010100;
				18'b011000011110001110: oled_data = 16'b1101110010110101;
				18'b011000100000001110: oled_data = 16'b1101110011010110;
				18'b011000100010001110: oled_data = 16'b1101110011010110;
				18'b011000100100001110: oled_data = 16'b1101110010010101;
				18'b011000100110001110: oled_data = 16'b1101010010010101;
				18'b011000101000001110: oled_data = 16'b1101110011010110;
				18'b011000101010001110: oled_data = 16'b1101110011010101;
				18'b011000101100001110: oled_data = 16'b1101110011010110;
				18'b011000101110001110: oled_data = 16'b1101110010110101;
				18'b011000110000001110: oled_data = 16'b1101110010010101;
				18'b011000110010001110: oled_data = 16'b1101110011010101;
				18'b011000110100001110: oled_data = 16'b1101110011010101;
				18'b011000110110001110: oled_data = 16'b1101110011010101;
				18'b011000111000001110: oled_data = 16'b1101110011010101;
				18'b011000111010001110: oled_data = 16'b1101110011010101;
				18'b011000111100001110: oled_data = 16'b1101110011010101;
				18'b011000111110001110: oled_data = 16'b1101110011010101;
				18'b011001000000001110: oled_data = 16'b1101110011010101;
				18'b011001000010001110: oled_data = 16'b1101010010010100;
				18'b011001000100001110: oled_data = 16'b1101110011010110;
				18'b011001000110001110: oled_data = 16'b1101110011010101;
				18'b011001001000001110: oled_data = 16'b1101110011010101;
				18'b011001001010001110: oled_data = 16'b1101110011010101;
				18'b011001001100001110: oled_data = 16'b1101110011010101;
				18'b011001001110001110: oled_data = 16'b1101110011010101;
				18'b011001010000001110: oled_data = 16'b1101110011010101;
				18'b011001010010001110: oled_data = 16'b1101110011010101;
				18'b011001010100001110: oled_data = 16'b1101110011010101;
				18'b011001010110001110: oled_data = 16'b1101110011010101;
				18'b011001011000001110: oled_data = 16'b1101110011010101;
				18'b011001011010001110: oled_data = 16'b1101110011010101;
				18'b011001011100001110: oled_data = 16'b1101110011010101;
				18'b011001011110001110: oled_data = 16'b1101110011010101;
				18'b011001100000001110: oled_data = 16'b1101110011010101;
				18'b011001100010001110: oled_data = 16'b1101110011010101;
				18'b011001100100001110: oled_data = 16'b1101110011010101;
				18'b011001100110001110: oled_data = 16'b1101110011010101;
				18'b011001101000001110: oled_data = 16'b1101110011010101;
				18'b011001101010001110: oled_data = 16'b1101110011010101;
				18'b011001101100001110: oled_data = 16'b1101110011010101;
				18'b011001101110001110: oled_data = 16'b1101110011010110;
				18'b011001110000001110: oled_data = 16'b1101110011010110;
				18'b011001110010001110: oled_data = 16'b1110010011010110;
				18'b011001110100001110: oled_data = 16'b1110010011010110;
				18'b011001110110001110: oled_data = 16'b1110010011010110;
				18'b011001111000001110: oled_data = 16'b1101110011010110;
				18'b011001111010001110: oled_data = 16'b1110010100010110;
				18'b011001111100001110: oled_data = 16'b1101110111011000;
				18'b011001111110001110: oled_data = 16'b0101101010101001;
				18'b011010000000001110: oled_data = 16'b0011100111000101;
				18'b011010000010001110: oled_data = 16'b0011000110000101;
				18'b011010000100001110: oled_data = 16'b0010100101000100;
				18'b011010000110001110: oled_data = 16'b0010000100000100;
				18'b011010001000001110: oled_data = 16'b0001100011100100;
				18'b011010001010001110: oled_data = 16'b0001100011100100;
				18'b011010001100001110: oled_data = 16'b0001100100100100;
				18'b011010001110001110: oled_data = 16'b0010000100100101;
				18'b011010010000001110: oled_data = 16'b0010000101000110;
				18'b011010010010001110: oled_data = 16'b0010000100100101;
				18'b011010010100001110: oled_data = 16'b0110001001101010;
				18'b011010010110001110: oled_data = 16'b1101010010010010;
				18'b011010011000001110: oled_data = 16'b1110110011110100;
				18'b011010011010001110: oled_data = 16'b1101001111001111;
				18'b011010011100001110: oled_data = 16'b1011101010001010;
				18'b011010011110001110: oled_data = 16'b1011001000001000;
				18'b011010100000001110: oled_data = 16'b1011001000101001;
				18'b011010100010001110: oled_data = 16'b1011001000101000;
				18'b011010100100001110: oled_data = 16'b1010101000101000;
				18'b011010100110001110: oled_data = 16'b1010101000001000;
				18'b011000011000001111: oled_data = 16'b1010111011111011;
				18'b011000011010001111: oled_data = 16'b1011110110011000;
				18'b011000011100001111: oled_data = 16'b1101010001010100;
				18'b011000011110001111: oled_data = 16'b1101110011010101;
				18'b011000100000001111: oled_data = 16'b1101110011010101;
				18'b011000100010001111: oled_data = 16'b1101110011010110;
				18'b011000100100001111: oled_data = 16'b1101010001110100;
				18'b011000100110001111: oled_data = 16'b1101110010110101;
				18'b011000101000001111: oled_data = 16'b1101110011010101;
				18'b011000101010001111: oled_data = 16'b1101110011010101;
				18'b011000101100001111: oled_data = 16'b1101110011010110;
				18'b011000101110001111: oled_data = 16'b1101010001010100;
				18'b011000110000001111: oled_data = 16'b1101110011010101;
				18'b011000110010001111: oled_data = 16'b1101110011010101;
				18'b011000110100001111: oled_data = 16'b1101110011010101;
				18'b011000110110001111: oled_data = 16'b1101110011010101;
				18'b011000111000001111: oled_data = 16'b1101110011010101;
				18'b011000111010001111: oled_data = 16'b1101110011010101;
				18'b011000111100001111: oled_data = 16'b1101110011010101;
				18'b011000111110001111: oled_data = 16'b1101110011010101;
				18'b011001000000001111: oled_data = 16'b1101110011010110;
				18'b011001000010001111: oled_data = 16'b1101010001110100;
				18'b011001000100001111: oled_data = 16'b1101110010110101;
				18'b011001000110001111: oled_data = 16'b1101110011010110;
				18'b011001001000001111: oled_data = 16'b1101110011010101;
				18'b011001001010001111: oled_data = 16'b1101110011010101;
				18'b011001001100001111: oled_data = 16'b1101110011010101;
				18'b011001001110001111: oled_data = 16'b1101110011010101;
				18'b011001010000001111: oled_data = 16'b1101110011010101;
				18'b011001010010001111: oled_data = 16'b1101110011010101;
				18'b011001010100001111: oled_data = 16'b1101110011010101;
				18'b011001010110001111: oled_data = 16'b1101110011010101;
				18'b011001011000001111: oled_data = 16'b1101110011010101;
				18'b011001011010001111: oled_data = 16'b1101110011010101;
				18'b011001011100001111: oled_data = 16'b1101110011010101;
				18'b011001011110001111: oled_data = 16'b1110010011110110;
				18'b011001100000001111: oled_data = 16'b1110010011110110;
				18'b011001100010001111: oled_data = 16'b1101110011010101;
				18'b011001100100001111: oled_data = 16'b1101110011010101;
				18'b011001100110001111: oled_data = 16'b1101110011010101;
				18'b011001101000001111: oled_data = 16'b1101110011010101;
				18'b011001101010001111: oled_data = 16'b1101110011010101;
				18'b011001101100001111: oled_data = 16'b1101110011010101;
				18'b011001101110001111: oled_data = 16'b1101110011010110;
				18'b011001110000001111: oled_data = 16'b1101110011010110;
				18'b011001110010001111: oled_data = 16'b1110010011010110;
				18'b011001110100001111: oled_data = 16'b1110010011010110;
				18'b011001110110001111: oled_data = 16'b1110010011010110;
				18'b011001111000001111: oled_data = 16'b1110010011010110;
				18'b011001111010001111: oled_data = 16'b1101110011010110;
				18'b011001111100001111: oled_data = 16'b1110110110011000;
				18'b011001111110001111: oled_data = 16'b1010010001010001;
				18'b011010000000001111: oled_data = 16'b0010100100000100;
				18'b011010000010001111: oled_data = 16'b0010100100100101;
				18'b011010000100001111: oled_data = 16'b0010000100100100;
				18'b011010000110001111: oled_data = 16'b0010000100100100;
				18'b011010001000001111: oled_data = 16'b0001100011100100;
				18'b011010001010001111: oled_data = 16'b0001100011100100;
				18'b011010001100001111: oled_data = 16'b0001100100000100;
				18'b011010001110001111: oled_data = 16'b0001100100100101;
				18'b011010010000001111: oled_data = 16'b0001100100100101;
				18'b011010010010001111: oled_data = 16'b0111101100001100;
				18'b011010010100001111: oled_data = 16'b1110010100010100;
				18'b011010010110001111: oled_data = 16'b1110010010010010;
				18'b011010011000001111: oled_data = 16'b1100001100001100;
				18'b011010011010001111: oled_data = 16'b1011001000101001;
				18'b011010011100001111: oled_data = 16'b1011001000101001;
				18'b011010011110001111: oled_data = 16'b1011001000101001;
				18'b011010100000001111: oled_data = 16'b1011001000101001;
				18'b011010100010001111: oled_data = 16'b1011001000101000;
				18'b011010100100001111: oled_data = 16'b1010101000001000;
				18'b011010100110001111: oled_data = 16'b1010101000001000;
				18'b011000011000010000: oled_data = 16'b1011011011111011;
				18'b011000011010010000: oled_data = 16'b1100010011110110;
				18'b011000011100010000: oled_data = 16'b1101110010010101;
				18'b011000011110010000: oled_data = 16'b1101110011010110;
				18'b011000100000010000: oled_data = 16'b1101110011010110;
				18'b011000100010010000: oled_data = 16'b1101110011010110;
				18'b011000100100010000: oled_data = 16'b1101010001110100;
				18'b011000100110010000: oled_data = 16'b1101110011010101;
				18'b011000101000010000: oled_data = 16'b1101110011010101;
				18'b011000101010010000: oled_data = 16'b1101110011010101;
				18'b011000101100010000: oled_data = 16'b1101110010110101;
				18'b011000101110010000: oled_data = 16'b1100110000110011;
				18'b011000110000010000: oled_data = 16'b1101110011010110;
				18'b011000110010010000: oled_data = 16'b1101110011010101;
				18'b011000110100010000: oled_data = 16'b1101110011010101;
				18'b011000110110010000: oled_data = 16'b1101110011010101;
				18'b011000111000010000: oled_data = 16'b1101110011010101;
				18'b011000111010010000: oled_data = 16'b1101110011010101;
				18'b011000111100010000: oled_data = 16'b1101110011010101;
				18'b011000111110010000: oled_data = 16'b1101110011010101;
				18'b011001000000010000: oled_data = 16'b1101110011010101;
				18'b011001000010010000: oled_data = 16'b1101110010110101;
				18'b011001000100010000: oled_data = 16'b1101010010010100;
				18'b011001000110010000: oled_data = 16'b1101110011010110;
				18'b011001001000010000: oled_data = 16'b1101110011010101;
				18'b011001001010010000: oled_data = 16'b1101110011010110;
				18'b011001001100010000: oled_data = 16'b1101110011010110;
				18'b011001001110010000: oled_data = 16'b1101110011010101;
				18'b011001010000010000: oled_data = 16'b1101110011010101;
				18'b011001010010010000: oled_data = 16'b1101110011010101;
				18'b011001010100010000: oled_data = 16'b1101110011010101;
				18'b011001010110010000: oled_data = 16'b1101110011010101;
				18'b011001011000010000: oled_data = 16'b1101110011010101;
				18'b011001011010010000: oled_data = 16'b1101110011010101;
				18'b011001011100010000: oled_data = 16'b1101110011010101;
				18'b011001011110010000: oled_data = 16'b1101110011010110;
				18'b011001100000010000: oled_data = 16'b1110010011110110;
				18'b011001100010010000: oled_data = 16'b1101110011010101;
				18'b011001100100010000: oled_data = 16'b1101110011010101;
				18'b011001100110010000: oled_data = 16'b1101110011010101;
				18'b011001101000010000: oled_data = 16'b1101110011010101;
				18'b011001101010010000: oled_data = 16'b1101110011010101;
				18'b011001101100010000: oled_data = 16'b1101110011010101;
				18'b011001101110010000: oled_data = 16'b1101110011010110;
				18'b011001110000010000: oled_data = 16'b1101110011010110;
				18'b011001110010010000: oled_data = 16'b1101110011010110;
				18'b011001110100010000: oled_data = 16'b1101110011010110;
				18'b011001110110010000: oled_data = 16'b1101110011010110;
				18'b011001111000010000: oled_data = 16'b1101110011010110;
				18'b011001111010010000: oled_data = 16'b1101110011010110;
				18'b011001111100010000: oled_data = 16'b1110010011010110;
				18'b011001111110010000: oled_data = 16'b1110010110010111;
				18'b011010000000010000: oled_data = 16'b0100101000001000;
				18'b011010000010010000: oled_data = 16'b0010000100100100;
				18'b011010000100010000: oled_data = 16'b0010100101100101;
				18'b011010000110010000: oled_data = 16'b0010100101100101;
				18'b011010001000010000: oled_data = 16'b0010000100000100;
				18'b011010001010010000: oled_data = 16'b0001100011100100;
				18'b011010001100010000: oled_data = 16'b0010000100100101;
				18'b011010001110010000: oled_data = 16'b0010000100100101;
				18'b011010010000010000: oled_data = 16'b1000101101001101;
				18'b011010010010010000: oled_data = 16'b1110110100110101;
				18'b011010010100010000: oled_data = 16'b1101110001010001;
				18'b011010010110010000: oled_data = 16'b1011101010101010;
				18'b011010011000010000: oled_data = 16'b1011001000101001;
				18'b011010011010010000: oled_data = 16'b1011001000101001;
				18'b011010011100010000: oled_data = 16'b1011001001001001;
				18'b011010011110010000: oled_data = 16'b1011001000101001;
				18'b011010100000010000: oled_data = 16'b1011001000101001;
				18'b011010100010010000: oled_data = 16'b1011001000101000;
				18'b011010100100010000: oled_data = 16'b1010101000001000;
				18'b011010100110010000: oled_data = 16'b1010101000001000;
				18'b011000011000010001: oled_data = 16'b1000110101010110;
				18'b011000011010010001: oled_data = 16'b1100010001110100;
				18'b011000011100010001: oled_data = 16'b1101110010110101;
				18'b011000011110010001: oled_data = 16'b1101110011010110;
				18'b011000100000010001: oled_data = 16'b1101110011010110;
				18'b011000100010010001: oled_data = 16'b1101110011010101;
				18'b011000100100010001: oled_data = 16'b1101010001110100;
				18'b011000100110010001: oled_data = 16'b1101110011010101;
				18'b011000101000010001: oled_data = 16'b1110010011110110;
				18'b011000101010010001: oled_data = 16'b1101110011010110;
				18'b011000101100010001: oled_data = 16'b1101010010010100;
				18'b011000101110010001: oled_data = 16'b1101010001110100;
				18'b011000110000010001: oled_data = 16'b1101110011010110;
				18'b011000110010010001: oled_data = 16'b1101110011010101;
				18'b011000110100010001: oled_data = 16'b1101110011010101;
				18'b011000110110010001: oled_data = 16'b1101110011010101;
				18'b011000111000010001: oled_data = 16'b1101110011010101;
				18'b011000111010010001: oled_data = 16'b1101110011010101;
				18'b011000111100010001: oled_data = 16'b1101110011010101;
				18'b011000111110010001: oled_data = 16'b1101110011010101;
				18'b011001000000010001: oled_data = 16'b1101110011010101;
				18'b011001000010010001: oled_data = 16'b1101110011010110;
				18'b011001000100010001: oled_data = 16'b1101010010010100;
				18'b011001000110010001: oled_data = 16'b1101110010110101;
				18'b011001001000010001: oled_data = 16'b1101110011010101;
				18'b011001001010010001: oled_data = 16'b1110010011010110;
				18'b011001001100010001: oled_data = 16'b1110010011010110;
				18'b011001001110010001: oled_data = 16'b1101110011010101;
				18'b011001010000010001: oled_data = 16'b1101110011010101;
				18'b011001010010010001: oled_data = 16'b1101110011010101;
				18'b011001010100010001: oled_data = 16'b1101110011010101;
				18'b011001010110010001: oled_data = 16'b1101110011010110;
				18'b011001011000010001: oled_data = 16'b1101110011010110;
				18'b011001011010010001: oled_data = 16'b1101110011010101;
				18'b011001011100010001: oled_data = 16'b1101110011010101;
				18'b011001011110010001: oled_data = 16'b1101110011010101;
				18'b011001100000010001: oled_data = 16'b1101110011010101;
				18'b011001100010010001: oled_data = 16'b1101110011010101;
				18'b011001100100010001: oled_data = 16'b1101110011010101;
				18'b011001100110010001: oled_data = 16'b1101110011010101;
				18'b011001101000010001: oled_data = 16'b1101110011010101;
				18'b011001101010010001: oled_data = 16'b1101110011010101;
				18'b011001101100010001: oled_data = 16'b1101110011010101;
				18'b011001101110010001: oled_data = 16'b1101110011010101;
				18'b011001110000010001: oled_data = 16'b1101110011010101;
				18'b011001110010010001: oled_data = 16'b1101110011010101;
				18'b011001110100010001: oled_data = 16'b1101110011010101;
				18'b011001110110010001: oled_data = 16'b1101110011010101;
				18'b011001111000010001: oled_data = 16'b1101110011010110;
				18'b011001111010010001: oled_data = 16'b1101110011010110;
				18'b011001111100010001: oled_data = 16'b1101110011010101;
				18'b011001111110010001: oled_data = 16'b1110110101010111;
				18'b011010000000010001: oled_data = 16'b1010010000010001;
				18'b011010000010010001: oled_data = 16'b0010100101000101;
				18'b011010000100010001: oled_data = 16'b0010100101100110;
				18'b011010000110010001: oled_data = 16'b0011000110000110;
				18'b011010001000010001: oled_data = 16'b0010100101000101;
				18'b011010001010010001: oled_data = 16'b0010000100000100;
				18'b011010001100010001: oled_data = 16'b0010000100100100;
				18'b011010001110010001: oled_data = 16'b1000101100101101;
				18'b011010010000010001: oled_data = 16'b1110110100010101;
				18'b011010010010010001: oled_data = 16'b1101110000010000;
				18'b011010010100010001: oled_data = 16'b1011001001101010;
				18'b011010010110010001: oled_data = 16'b1011001001001001;
				18'b011010011000010001: oled_data = 16'b1011001001001001;
				18'b011010011010010001: oled_data = 16'b1011001000101001;
				18'b011010011100010001: oled_data = 16'b1011001000101001;
				18'b011010011110010001: oled_data = 16'b1011001000101001;
				18'b011010100000010001: oled_data = 16'b1011001000101001;
				18'b011010100010010001: oled_data = 16'b1011001000101000;
				18'b011010100100010001: oled_data = 16'b1011001000001000;
				18'b011010100110010001: oled_data = 16'b1011001000001000;
				18'b011000011000010010: oled_data = 16'b0111010001010011;
				18'b011000011010010010: oled_data = 16'b1101010010010100;
				18'b011000011100010010: oled_data = 16'b1101110011010101;
				18'b011000011110010010: oled_data = 16'b1101110011010110;
				18'b011000100000010010: oled_data = 16'b1101110011010110;
				18'b011000100010010010: oled_data = 16'b1101110010110101;
				18'b011000100100010010: oled_data = 16'b1101010010010101;
				18'b011000100110010010: oled_data = 16'b1110010011010110;
				18'b011000101000010010: oled_data = 16'b1110010100010110;
				18'b011000101010010010: oled_data = 16'b1101110011010110;
				18'b011000101100010010: oled_data = 16'b1101010001110100;
				18'b011000101110010010: oled_data = 16'b1101110010010101;
				18'b011000110000010010: oled_data = 16'b1101110011010110;
				18'b011000110010010010: oled_data = 16'b1101110011010101;
				18'b011000110100010010: oled_data = 16'b1101110011010101;
				18'b011000110110010010: oled_data = 16'b1101110011010101;
				18'b011000111000010010: oled_data = 16'b1101110011010101;
				18'b011000111010010010: oled_data = 16'b1101110011010101;
				18'b011000111100010010: oled_data = 16'b1101110011010101;
				18'b011000111110010010: oled_data = 16'b1101110011010101;
				18'b011001000000010010: oled_data = 16'b1101110011010101;
				18'b011001000010010010: oled_data = 16'b1101110011010110;
				18'b011001000100010010: oled_data = 16'b1101110010010101;
				18'b011001000110010010: oled_data = 16'b1101010001110100;
				18'b011001001000010010: oled_data = 16'b1101110011010110;
				18'b011001001010010010: oled_data = 16'b1101110011010110;
				18'b011001001100010010: oled_data = 16'b1101110011010110;
				18'b011001001110010010: oled_data = 16'b1101110011010101;
				18'b011001010000010010: oled_data = 16'b1101110011010101;
				18'b011001010010010010: oled_data = 16'b1101110011010101;
				18'b011001010100010010: oled_data = 16'b1101110011010101;
				18'b011001010110010010: oled_data = 16'b1110010011110110;
				18'b011001011000010010: oled_data = 16'b1110110100110111;
				18'b011001011010010010: oled_data = 16'b1101110011010110;
				18'b011001011100010010: oled_data = 16'b1101110011010101;
				18'b011001011110010010: oled_data = 16'b1101110011010101;
				18'b011001100000010010: oled_data = 16'b1101110011010101;
				18'b011001100010010010: oled_data = 16'b1101110011010101;
				18'b011001100100010010: oled_data = 16'b1101110011010101;
				18'b011001100110010010: oled_data = 16'b1101110011010101;
				18'b011001101000010010: oled_data = 16'b1101110011010101;
				18'b011001101010010010: oled_data = 16'b1101110011010101;
				18'b011001101100010010: oled_data = 16'b1101110011010101;
				18'b011001101110010010: oled_data = 16'b1101110011010101;
				18'b011001110000010010: oled_data = 16'b1101110011010101;
				18'b011001110010010010: oled_data = 16'b1101110011010101;
				18'b011001110100010010: oled_data = 16'b1101110011010101;
				18'b011001110110010010: oled_data = 16'b1101110011010110;
				18'b011001111000010010: oled_data = 16'b1101110011010110;
				18'b011001111010010010: oled_data = 16'b1101110011010110;
				18'b011001111100010010: oled_data = 16'b1101110011010110;
				18'b011001111110010010: oled_data = 16'b1101110011010110;
				18'b011010000000010010: oled_data = 16'b1101110101010111;
				18'b011010000010010010: oled_data = 16'b0101101000001001;
				18'b011010000100010010: oled_data = 16'b0010100101100110;
				18'b011010000110010010: oled_data = 16'b0011000110000110;
				18'b011010001000010010: oled_data = 16'b0010100101000101;
				18'b011010001010010010: oled_data = 16'b0010000100000100;
				18'b011010001100010010: oled_data = 16'b1000001100001101;
				18'b011010001110010010: oled_data = 16'b1110110100010100;
				18'b011010010000010010: oled_data = 16'b1101110000010000;
				18'b011010010010010010: oled_data = 16'b1011001001101001;
				18'b011010010100010010: oled_data = 16'b1011001001001001;
				18'b011010010110010010: oled_data = 16'b1011001001001001;
				18'b011010011000010010: oled_data = 16'b1011001001001001;
				18'b011010011010010010: oled_data = 16'b1011001000101001;
				18'b011010011100010010: oled_data = 16'b1011001000101001;
				18'b011010011110010010: oled_data = 16'b1011001000101001;
				18'b011010100000010010: oled_data = 16'b1011001000101001;
				18'b011010100010010010: oled_data = 16'b1011001000101000;
				18'b011010100100010010: oled_data = 16'b1011001000101000;
				18'b011010100110010010: oled_data = 16'b1011001000001000;
				18'b011000011000010011: oled_data = 16'b1001010000110100;
				18'b011000011010010011: oled_data = 16'b1101110010110101;
				18'b011000011100010011: oled_data = 16'b1101110011010110;
				18'b011000011110010011: oled_data = 16'b1101110011010101;
				18'b011000100000010011: oled_data = 16'b1101110011010101;
				18'b011000100010010011: oled_data = 16'b1101010010010101;
				18'b011000100100010011: oled_data = 16'b1101010010010100;
				18'b011000100110010011: oled_data = 16'b1110010011110110;
				18'b011000101000010011: oled_data = 16'b1110010011110110;
				18'b011000101010010011: oled_data = 16'b1101110011010101;
				18'b011000101100010011: oled_data = 16'b1100110001010011;
				18'b011000101110010011: oled_data = 16'b1101110010110101;
				18'b011000110000010011: oled_data = 16'b1101110011010101;
				18'b011000110010010011: oled_data = 16'b1101110011010101;
				18'b011000110100010011: oled_data = 16'b1101110011010101;
				18'b011000110110010011: oled_data = 16'b1110010100010110;
				18'b011000111000010011: oled_data = 16'b1101110011010110;
				18'b011000111010010011: oled_data = 16'b1101110011010101;
				18'b011000111100010011: oled_data = 16'b1101110011010101;
				18'b011000111110010011: oled_data = 16'b1101110011010101;
				18'b011001000000010011: oled_data = 16'b1101110011010101;
				18'b011001000010010011: oled_data = 16'b1101110011010101;
				18'b011001000100010011: oled_data = 16'b1101110011010110;
				18'b011001000110010011: oled_data = 16'b1100110001010011;
				18'b011001001000010011: oled_data = 16'b1101110011010101;
				18'b011001001010010011: oled_data = 16'b1101110011010101;
				18'b011001001100010011: oled_data = 16'b1101110011010101;
				18'b011001001110010011: oled_data = 16'b1101110011010101;
				18'b011001010000010011: oled_data = 16'b1101110011010101;
				18'b011001010010010011: oled_data = 16'b1101110010110101;
				18'b011001010100010011: oled_data = 16'b1101110011010101;
				18'b011001010110010011: oled_data = 16'b1101110011010101;
				18'b011001011000010011: oled_data = 16'b1110010011110110;
				18'b011001011010010011: oled_data = 16'b1101110011010110;
				18'b011001011100010011: oled_data = 16'b1101110011010110;
				18'b011001011110010011: oled_data = 16'b1101110011010101;
				18'b011001100000010011: oled_data = 16'b1101110011010101;
				18'b011001100010010011: oled_data = 16'b1101110011010101;
				18'b011001100100010011: oled_data = 16'b1101110011010101;
				18'b011001100110010011: oled_data = 16'b1101110011010101;
				18'b011001101000010011: oled_data = 16'b1101110011010101;
				18'b011001101010010011: oled_data = 16'b1101110011010101;
				18'b011001101100010011: oled_data = 16'b1101110011010101;
				18'b011001101110010011: oled_data = 16'b1101110011010101;
				18'b011001110000010011: oled_data = 16'b1101110011010101;
				18'b011001110010010011: oled_data = 16'b1101110011010110;
				18'b011001110100010011: oled_data = 16'b1101110011010101;
				18'b011001110110010011: oled_data = 16'b1101110011010110;
				18'b011001111000010011: oled_data = 16'b1101110011010101;
				18'b011001111010010011: oled_data = 16'b1101110011010101;
				18'b011001111100010011: oled_data = 16'b1101110011010101;
				18'b011001111110010011: oled_data = 16'b1101110011010101;
				18'b011010000000010011: oled_data = 16'b1110010011110110;
				18'b011010000010010011: oled_data = 16'b1010001111010000;
				18'b011010000100010011: oled_data = 16'b0011000101100101;
				18'b011010000110010011: oled_data = 16'b0011000110000110;
				18'b011010001000010011: oled_data = 16'b0010000100000100;
				18'b011010001010010011: oled_data = 16'b0110001010001010;
				18'b011010001100010011: oled_data = 16'b1110010100010101;
				18'b011010001110010011: oled_data = 16'b1110010001010001;
				18'b011010010000010011: oled_data = 16'b1011001010001010;
				18'b011010010010010011: oled_data = 16'b1011001001001001;
				18'b011010010100010011: oled_data = 16'b1011001001001001;
				18'b011010010110010011: oled_data = 16'b1011001001001001;
				18'b011010011000010011: oled_data = 16'b1011001001001001;
				18'b011010011010010011: oled_data = 16'b1011001000101001;
				18'b011010011100010011: oled_data = 16'b1011001000101001;
				18'b011010011110010011: oled_data = 16'b1011001000101001;
				18'b011010100000010011: oled_data = 16'b1011001000101001;
				18'b011010100010010011: oled_data = 16'b1011001000101001;
				18'b011010100100010011: oled_data = 16'b1011001000101000;
				18'b011010100110010011: oled_data = 16'b1011001000001000;
				18'b011000011000010100: oled_data = 16'b1011010001010100;
				18'b011000011010010100: oled_data = 16'b1110010010110101;
				18'b011000011100010100: oled_data = 16'b1101110010110101;
				18'b011000011110010100: oled_data = 16'b1101110010110101;
				18'b011000100000010100: oled_data = 16'b1101110011010110;
				18'b011000100010010100: oled_data = 16'b1100110001010011;
				18'b011000100100010100: oled_data = 16'b1101010001110100;
				18'b011000100110010100: oled_data = 16'b1110010011110110;
				18'b011000101000010100: oled_data = 16'b1110010011110110;
				18'b011000101010010100: oled_data = 16'b1101110011010101;
				18'b011000101100010100: oled_data = 16'b1100110001010011;
				18'b011000101110010100: oled_data = 16'b1101110010110101;
				18'b011000110000010100: oled_data = 16'b1101110011010101;
				18'b011000110010010100: oled_data = 16'b1101110011010101;
				18'b011000110100010100: oled_data = 16'b1101110011010101;
				18'b011000110110010100: oled_data = 16'b1110110110011000;
				18'b011000111000010100: oled_data = 16'b1110010100010110;
				18'b011000111010010100: oled_data = 16'b1101110011010101;
				18'b011000111100010100: oled_data = 16'b1101110011010101;
				18'b011000111110010100: oled_data = 16'b1101110011010101;
				18'b011001000000010100: oled_data = 16'b1101110011010101;
				18'b011001000010010100: oled_data = 16'b1101110011010101;
				18'b011001000100010100: oled_data = 16'b1110010011010110;
				18'b011001000110010100: oled_data = 16'b1100110001010011;
				18'b011001001000010100: oled_data = 16'b1101010001110100;
				18'b011001001010010100: oled_data = 16'b1101110011010110;
				18'b011001001100010100: oled_data = 16'b1101110011010101;
				18'b011001001110010100: oled_data = 16'b1101110011010101;
				18'b011001010000010100: oled_data = 16'b1101110011010101;
				18'b011001010010010100: oled_data = 16'b1101010010010100;
				18'b011001010100010100: oled_data = 16'b1101110011010101;
				18'b011001010110010100: oled_data = 16'b1101110011010101;
				18'b011001011000010100: oled_data = 16'b1101110011010101;
				18'b011001011010010100: oled_data = 16'b1101110011010101;
				18'b011001011100010100: oled_data = 16'b1101110011010101;
				18'b011001011110010100: oled_data = 16'b1101110011010101;
				18'b011001100000010100: oled_data = 16'b1101110011010110;
				18'b011001100010010100: oled_data = 16'b1101110011010101;
				18'b011001100100010100: oled_data = 16'b1101110011010101;
				18'b011001100110010100: oled_data = 16'b1101110011010101;
				18'b011001101000010100: oled_data = 16'b1101110011010101;
				18'b011001101010010100: oled_data = 16'b1101110011010101;
				18'b011001101100010100: oled_data = 16'b1101110011010101;
				18'b011001101110010100: oled_data = 16'b1101110011010101;
				18'b011001110000010100: oled_data = 16'b1101110011010101;
				18'b011001110010010100: oled_data = 16'b1101110011010101;
				18'b011001110100010100: oled_data = 16'b1101110011010101;
				18'b011001110110010100: oled_data = 16'b1101110011010101;
				18'b011001111000010100: oled_data = 16'b1101110011010110;
				18'b011001111010010100: oled_data = 16'b1101110010110101;
				18'b011001111100010100: oled_data = 16'b1101110010110101;
				18'b011001111110010100: oled_data = 16'b1101110011010110;
				18'b011010000000010100: oled_data = 16'b1110010011010110;
				18'b011010000010010100: oled_data = 16'b1101110011110110;
				18'b011010000100010100: oled_data = 16'b0110001010101011;
				18'b011010000110010100: oled_data = 16'b0010000100100101;
				18'b011010001000010100: oled_data = 16'b0101001000001000;
				18'b011010001010010100: oled_data = 16'b1101110011010100;
				18'b011010001100010100: oled_data = 16'b1110010010010010;
				18'b011010001110010100: oled_data = 16'b1011101010101011;
				18'b011010010000010100: oled_data = 16'b1011001001001001;
				18'b011010010010010100: oled_data = 16'b1011001001001001;
				18'b011010010100010100: oled_data = 16'b1011001001001001;
				18'b011010010110010100: oled_data = 16'b1011001001001001;
				18'b011010011000010100: oled_data = 16'b1011001001001001;
				18'b011010011010010100: oled_data = 16'b1011001000101001;
				18'b011010011100010100: oled_data = 16'b1011001000101001;
				18'b011010011110010100: oled_data = 16'b1011001000101001;
				18'b011010100000010100: oled_data = 16'b1010101000101000;
				18'b011010100010010100: oled_data = 16'b1011001000101001;
				18'b011010100100010100: oled_data = 16'b1011001000101000;
				18'b011010100110010100: oled_data = 16'b1011001000001000;
				18'b011000011000010101: oled_data = 16'b1011110001010100;
				18'b011000011010010101: oled_data = 16'b1101110011010101;
				18'b011000011100010101: oled_data = 16'b1101010010010100;
				18'b011000011110010101: oled_data = 16'b1101110011010110;
				18'b011000100000010101: oled_data = 16'b1110010011010110;
				18'b011000100010010101: oled_data = 16'b1100110000110011;
				18'b011000100100010101: oled_data = 16'b1101010010010101;
				18'b011000100110010101: oled_data = 16'b1101110011010110;
				18'b011000101000010101: oled_data = 16'b1101110011010101;
				18'b011000101010010101: oled_data = 16'b1101010011010100;
				18'b011000101100010101: oled_data = 16'b1100010001110010;
				18'b011000101110010101: oled_data = 16'b1101110010110101;
				18'b011000110000010101: oled_data = 16'b1101110011010101;
				18'b011000110010010101: oled_data = 16'b1101110011010101;
				18'b011000110100010101: oled_data = 16'b1101110011010101;
				18'b011000110110010101: oled_data = 16'b1110010101010111;
				18'b011000111000010101: oled_data = 16'b1110010100010110;
				18'b011000111010010101: oled_data = 16'b1101110011010101;
				18'b011000111100010101: oled_data = 16'b1101110011010101;
				18'b011000111110010101: oled_data = 16'b1101110011010101;
				18'b011001000000010101: oled_data = 16'b1101110011010101;
				18'b011001000010010101: oled_data = 16'b1101110011010101;
				18'b011001000100010101: oled_data = 16'b1101110011010101;
				18'b011001000110010101: oled_data = 16'b1101110010110101;
				18'b011001001000010101: oled_data = 16'b1100110000110011;
				18'b011001001010010101: oled_data = 16'b1110010011010110;
				18'b011001001100010101: oled_data = 16'b1101110011010101;
				18'b011001001110010101: oled_data = 16'b1101110011010110;
				18'b011001010000010101: oled_data = 16'b1101110011010110;
				18'b011001010010010101: oled_data = 16'b1101110010110101;
				18'b011001010100010101: oled_data = 16'b1101110010110101;
				18'b011001010110010101: oled_data = 16'b1101110011010110;
				18'b011001011000010101: oled_data = 16'b1101110011010101;
				18'b011001011010010101: oled_data = 16'b1101110011010101;
				18'b011001011100010101: oled_data = 16'b1101110011010101;
				18'b011001011110010101: oled_data = 16'b1101110010010101;
				18'b011001100000010101: oled_data = 16'b1101110010010101;
				18'b011001100010010101: oled_data = 16'b1101110011010101;
				18'b011001100100010101: oled_data = 16'b1101110011010110;
				18'b011001100110010101: oled_data = 16'b1101110011010101;
				18'b011001101000010101: oled_data = 16'b1101110011010101;
				18'b011001101010010101: oled_data = 16'b1101110011010101;
				18'b011001101100010101: oled_data = 16'b1101110011010101;
				18'b011001101110010101: oled_data = 16'b1101110011010101;
				18'b011001110000010101: oled_data = 16'b1101110011010101;
				18'b011001110010010101: oled_data = 16'b1101110011010101;
				18'b011001110100010101: oled_data = 16'b1101110011010101;
				18'b011001110110010101: oled_data = 16'b1101110011010101;
				18'b011001111000010101: oled_data = 16'b1101110011010110;
				18'b011001111010010101: oled_data = 16'b1101110011010110;
				18'b011001111100010101: oled_data = 16'b1101010010010100;
				18'b011001111110010101: oled_data = 16'b1101010010010100;
				18'b011010000000010101: oled_data = 16'b1110010011010110;
				18'b011010000010010101: oled_data = 16'b1110010011010110;
				18'b011010000100010101: oled_data = 16'b1100110010010100;
				18'b011010000110010101: oled_data = 16'b0101100111101001;
				18'b011010001000010101: oled_data = 16'b1011010000110001;
				18'b011010001010010101: oled_data = 16'b1110110100010100;
				18'b011010001100010101: oled_data = 16'b1100001100101101;
				18'b011010001110010101: oled_data = 16'b1011001000101001;
				18'b011010010000010101: oled_data = 16'b1011101001001001;
				18'b011010010010010101: oled_data = 16'b1011101001001001;
				18'b011010010100010101: oled_data = 16'b1011001000101001;
				18'b011010010110010101: oled_data = 16'b1011001001001001;
				18'b011010011000010101: oled_data = 16'b1011001001001001;
				18'b011010011010010101: oled_data = 16'b1011001001001001;
				18'b011010011100010101: oled_data = 16'b1011001000101001;
				18'b011010011110010101: oled_data = 16'b1010001000001000;
				18'b011010100000010101: oled_data = 16'b1010101000101000;
				18'b011010100010010101: oled_data = 16'b1011001000101001;
				18'b011010100100010101: oled_data = 16'b1011001000101000;
				18'b011010100110010101: oled_data = 16'b1011001000001000;
				18'b011000011000010110: oled_data = 16'b1101010010010100;
				18'b011000011010010110: oled_data = 16'b1101110010110101;
				18'b011000011100010110: oled_data = 16'b1100110000110011;
				18'b011000011110010110: oled_data = 16'b1110010011110110;
				18'b011000100000010110: oled_data = 16'b1110010011010110;
				18'b011000100010010110: oled_data = 16'b1100010000010010;
				18'b011000100100010110: oled_data = 16'b1101010010010101;
				18'b011000100110010110: oled_data = 16'b1101110011010110;
				18'b011000101000010110: oled_data = 16'b1101110011010101;
				18'b011000101010010110: oled_data = 16'b1101010011010100;
				18'b011000101100010110: oled_data = 16'b1100110010110011;
				18'b011000101110010110: oled_data = 16'b1101110010110101;
				18'b011000110000010110: oled_data = 16'b1101110010110101;
				18'b011000110010010110: oled_data = 16'b1101110010110101;
				18'b011000110100010110: oled_data = 16'b1101110011010101;
				18'b011000110110010110: oled_data = 16'b1110010100010110;
				18'b011000111000010110: oled_data = 16'b1110010011110110;
				18'b011000111010010110: oled_data = 16'b1101110011010101;
				18'b011000111100010110: oled_data = 16'b1101110011010101;
				18'b011000111110010110: oled_data = 16'b1101110011010101;
				18'b011001000000010110: oled_data = 16'b1101110011010101;
				18'b011001000010010110: oled_data = 16'b1101110011010101;
				18'b011001000100010110: oled_data = 16'b1101110011010101;
				18'b011001000110010110: oled_data = 16'b1101110011010110;
				18'b011001001000010110: oled_data = 16'b1100001111110010;
				18'b011001001010010110: oled_data = 16'b1101110010110101;
				18'b011001001100010110: oled_data = 16'b1101110011010110;
				18'b011001001110010110: oled_data = 16'b1101110011010110;
				18'b011001010000010110: oled_data = 16'b1101110011010101;
				18'b011001010010010110: oled_data = 16'b1101110011010101;
				18'b011001010100010110: oled_data = 16'b1101010001110100;
				18'b011001010110010110: oled_data = 16'b1101110011010101;
				18'b011001011000010110: oled_data = 16'b1101110011010101;
				18'b011001011010010110: oled_data = 16'b1101110011010101;
				18'b011001011100010110: oled_data = 16'b1101110011010101;
				18'b011001011110010110: oled_data = 16'b1101110011010101;
				18'b011001100000010110: oled_data = 16'b1101010010010101;
				18'b011001100010010110: oled_data = 16'b1101010001110100;
				18'b011001100100010110: oled_data = 16'b1101010010010101;
				18'b011001100110010110: oled_data = 16'b1101110011010101;
				18'b011001101000010110: oled_data = 16'b1101110011010110;
				18'b011001101010010110: oled_data = 16'b1101110011010110;
				18'b011001101100010110: oled_data = 16'b1101110011010110;
				18'b011001101110010110: oled_data = 16'b1101110011010101;
				18'b011001110000010110: oled_data = 16'b1101110011010101;
				18'b011001110010010110: oled_data = 16'b1101110011010101;
				18'b011001110100010110: oled_data = 16'b1101110011010101;
				18'b011001110110010110: oled_data = 16'b1101110011010110;
				18'b011001111000010110: oled_data = 16'b1101110011010110;
				18'b011001111010010110: oled_data = 16'b1101110011010110;
				18'b011001111100010110: oled_data = 16'b1101110011010110;
				18'b011001111110010110: oled_data = 16'b1101010010010100;
				18'b011010000000010110: oled_data = 16'b1101010010010100;
				18'b011010000010010110: oled_data = 16'b1101110011010101;
				18'b011010000100010110: oled_data = 16'b1101110011010101;
				18'b011010000110010110: oled_data = 16'b1100110001110011;
				18'b011010001000010110: oled_data = 16'b1110110100010100;
				18'b011010001010010110: oled_data = 16'b1101001111101111;
				18'b011010001100010110: oled_data = 16'b1011001001001001;
				18'b011010001110010110: oled_data = 16'b1011101001001001;
				18'b011010010000010110: oled_data = 16'b1011101001001001;
				18'b011010010010010110: oled_data = 16'b1011101001001001;
				18'b011010010100010110: oled_data = 16'b1011001000101001;
				18'b011010010110010110: oled_data = 16'b1011001001001001;
				18'b011010011000010110: oled_data = 16'b1011001001001001;
				18'b011010011010010110: oled_data = 16'b1010101000101000;
				18'b011010011100010110: oled_data = 16'b1010001000001000;
				18'b011010011110010110: oled_data = 16'b1011001000101001;
				18'b011010100000010110: oled_data = 16'b1011001000101001;
				18'b011010100010010110: oled_data = 16'b1011001000101001;
				18'b011010100100010110: oled_data = 16'b1011001000101000;
				18'b011010100110010110: oled_data = 16'b1011001000001000;
				18'b011000011000010111: oled_data = 16'b1101010010010100;
				18'b011000011010010111: oled_data = 16'b1101110010110100;
				18'b011000011100010111: oled_data = 16'b1100110001110100;
				18'b011000011110010111: oled_data = 16'b1110010011110110;
				18'b011000100000010111: oled_data = 16'b1110010011010110;
				18'b011000100010010111: oled_data = 16'b1100110000010011;
				18'b011000100100010111: oled_data = 16'b1101110010110101;
				18'b011000100110010111: oled_data = 16'b1101110011010110;
				18'b011000101000010111: oled_data = 16'b1101110011010101;
				18'b011000101010010111: oled_data = 16'b1101110100010101;
				18'b011000101100010111: oled_data = 16'b1101010011110101;
				18'b011000101110010111: oled_data = 16'b1101110010110101;
				18'b011000110000010111: oled_data = 16'b1101110010110101;
				18'b011000110010010111: oled_data = 16'b1101010010010100;
				18'b011000110100010111: oled_data = 16'b1101110011010110;
				18'b011000110110010111: oled_data = 16'b1101110011010101;
				18'b011000111000010111: oled_data = 16'b1101110011010101;
				18'b011000111010010111: oled_data = 16'b1101110011010101;
				18'b011000111100010111: oled_data = 16'b1101110011010101;
				18'b011000111110010111: oled_data = 16'b1101110011010101;
				18'b011001000000010111: oled_data = 16'b1101110011010101;
				18'b011001000010010111: oled_data = 16'b1101010010010100;
				18'b011001000100010111: oled_data = 16'b1101110011010101;
				18'b011001000110010111: oled_data = 16'b1101110011010110;
				18'b011001001000010111: oled_data = 16'b1101010001110100;
				18'b011001001010010111: oled_data = 16'b1100110001010011;
				18'b011001001100010111: oled_data = 16'b1101110011110110;
				18'b011001001110010111: oled_data = 16'b1101110011010101;
				18'b011001010000010111: oled_data = 16'b1101110011010101;
				18'b011001010010010111: oled_data = 16'b1110010011010110;
				18'b011001010100010111: oled_data = 16'b1101010001010100;
				18'b011001010110010111: oled_data = 16'b1101010010110101;
				18'b011001011000010111: oled_data = 16'b1101110011010110;
				18'b011001011010010111: oled_data = 16'b1101110011010101;
				18'b011001011100010111: oled_data = 16'b1101110011010101;
				18'b011001011110010111: oled_data = 16'b1110010011010110;
				18'b011001100000010111: oled_data = 16'b1110010011110110;
				18'b011001100010010111: oled_data = 16'b1101110011010101;
				18'b011001100100010111: oled_data = 16'b1101010001110100;
				18'b011001100110010111: oled_data = 16'b1101010001110100;
				18'b011001101000010111: oled_data = 16'b1101010001110100;
				18'b011001101010010111: oled_data = 16'b1101010010010100;
				18'b011001101100010111: oled_data = 16'b1101110010110101;
				18'b011001101110010111: oled_data = 16'b1101110010110101;
				18'b011001110000010111: oled_data = 16'b1101110010110101;
				18'b011001110010010111: oled_data = 16'b1101110010110101;
				18'b011001110100010111: oled_data = 16'b1101110010010101;
				18'b011001110110010111: oled_data = 16'b1101010010010100;
				18'b011001111000010111: oled_data = 16'b1101110010110101;
				18'b011001111010010111: oled_data = 16'b1101110011010110;
				18'b011001111100010111: oled_data = 16'b1110010011010110;
				18'b011001111110010111: oled_data = 16'b1110010011010110;
				18'b011010000000010111: oled_data = 16'b1101110010110101;
				18'b011010000010010111: oled_data = 16'b1101010001110100;
				18'b011010000100010111: oled_data = 16'b1101010001110011;
				18'b011010000110010111: oled_data = 16'b1110010011110100;
				18'b011010001000010111: oled_data = 16'b1110010010110010;
				18'b011010001010010111: oled_data = 16'b1011101010001010;
				18'b011010001100010111: oled_data = 16'b1011001000101001;
				18'b011010001110010111: oled_data = 16'b1011001001001001;
				18'b011010010000010111: oled_data = 16'b1011001001001001;
				18'b011010010010010111: oled_data = 16'b1011001001001001;
				18'b011010010100010111: oled_data = 16'b1011001001001001;
				18'b011010010110010111: oled_data = 16'b1011001001001001;
				18'b011010011000010111: oled_data = 16'b1011001000101001;
				18'b011010011010010111: oled_data = 16'b1010101000001000;
				18'b011010011100010111: oled_data = 16'b1011001001001001;
				18'b011010011110010111: oled_data = 16'b1011001001001001;
				18'b011010100000010111: oled_data = 16'b1011001000101001;
				18'b011010100010010111: oled_data = 16'b1011001000101001;
				18'b011010100100010111: oled_data = 16'b1011001000101000;
				18'b011010100110010111: oled_data = 16'b1011001000001000;
				18'b011000011000011000: oled_data = 16'b1101110010110101;
				18'b011000011010011000: oled_data = 16'b1101010010110010;
				18'b011000011100011000: oled_data = 16'b1100110010010010;
				18'b011000011110011000: oled_data = 16'b1110010011010110;
				18'b011000100000011000: oled_data = 16'b1110010011010110;
				18'b011000100010011000: oled_data = 16'b1100110000010011;
				18'b011000100100011000: oled_data = 16'b1101110010110101;
				18'b011000100110011000: oled_data = 16'b1101110011010110;
				18'b011000101000011000: oled_data = 16'b1101110011010101;
				18'b011000101010011000: oled_data = 16'b1101010101010110;
				18'b011000101100011000: oled_data = 16'b1101010101110110;
				18'b011000101110011000: oled_data = 16'b1101110010010101;
				18'b011000110000011000: oled_data = 16'b1101110010110101;
				18'b011000110010011000: oled_data = 16'b1101010010010100;
				18'b011000110100011000: oled_data = 16'b1101110011010110;
				18'b011000110110011000: oled_data = 16'b1101110011010101;
				18'b011000111000011000: oled_data = 16'b1101110011010101;
				18'b011000111010011000: oled_data = 16'b1101110011010101;
				18'b011000111100011000: oled_data = 16'b1101110011010101;
				18'b011000111110011000: oled_data = 16'b1101110011010101;
				18'b011001000000011000: oled_data = 16'b1101110011110110;
				18'b011001000010011000: oled_data = 16'b1100110001010011;
				18'b011001000100011000: oled_data = 16'b1101010010010100;
				18'b011001000110011000: oled_data = 16'b1101110011010110;
				18'b011001001000011000: oled_data = 16'b1101110011010101;
				18'b011001001010011000: oled_data = 16'b1100010000010011;
				18'b011001001100011000: oled_data = 16'b1101110011010101;
				18'b011001001110011000: oled_data = 16'b1101110011010101;
				18'b011001010000011000: oled_data = 16'b1101110011010101;
				18'b011001010010011000: oled_data = 16'b1101110011010110;
				18'b011001010100011000: oled_data = 16'b1101010010010100;
				18'b011001010110011000: oled_data = 16'b1100110000110011;
				18'b011001011000011000: oled_data = 16'b1101110011010110;
				18'b011001011010011000: oled_data = 16'b1101110011010101;
				18'b011001011100011000: oled_data = 16'b1101110011010101;
				18'b011001011110011000: oled_data = 16'b1101110011010101;
				18'b011001100000011000: oled_data = 16'b1110010011010110;
				18'b011001100010011000: oled_data = 16'b1101110011010110;
				18'b011001100100011000: oled_data = 16'b1101110011010110;
				18'b011001100110011000: oled_data = 16'b1101110011010101;
				18'b011001101000011000: oled_data = 16'b1101110010110101;
				18'b011001101010011000: oled_data = 16'b1101010010010100;
				18'b011001101100011000: oled_data = 16'b1101010001110100;
				18'b011001101110011000: oled_data = 16'b1101010001110100;
				18'b011001110000011000: oled_data = 16'b1101010001010100;
				18'b011001110010011000: oled_data = 16'b1101010001010100;
				18'b011001110100011000: oled_data = 16'b1101010001110100;
				18'b011001110110011000: oled_data = 16'b1101010001010100;
				18'b011001111000011000: oled_data = 16'b1101110010110101;
				18'b011001111010011000: oled_data = 16'b1101110011010101;
				18'b011001111100011000: oled_data = 16'b1110010011010110;
				18'b011001111110011000: oled_data = 16'b1110010011010110;
				18'b011010000000011000: oled_data = 16'b1110010011110110;
				18'b011010000010011000: oled_data = 16'b1101110010010101;
				18'b011010000100011000: oled_data = 16'b1101010010010011;
				18'b011010000110011000: oled_data = 16'b1110110100010100;
				18'b011010001000011000: oled_data = 16'b1100101101101101;
				18'b011010001010011000: oled_data = 16'b1011001000101001;
				18'b011010001100011000: oled_data = 16'b1011001001001001;
				18'b011010001110011000: oled_data = 16'b1011001001001001;
				18'b011010010000011000: oled_data = 16'b1011001001001001;
				18'b011010010010011000: oled_data = 16'b1011001001001001;
				18'b011010010100011000: oled_data = 16'b1011001001001001;
				18'b011010010110011000: oled_data = 16'b1011001000101001;
				18'b011010011000011000: oled_data = 16'b1010101000001000;
				18'b011010011010011000: oled_data = 16'b1011001001001001;
				18'b011010011100011000: oled_data = 16'b1011001001001001;
				18'b011010011110011000: oled_data = 16'b1011001001001001;
				18'b011010100000011000: oled_data = 16'b1011001000101001;
				18'b011010100010011000: oled_data = 16'b1011001000101001;
				18'b011010100100011000: oled_data = 16'b1011001000101000;
				18'b011010100110011000: oled_data = 16'b1011001000001000;
				18'b011000011000011001: oled_data = 16'b1110010011110110;
				18'b011000011010011001: oled_data = 16'b1100010001010001;
				18'b011000011100011001: oled_data = 16'b1100110001110010;
				18'b011000011110011001: oled_data = 16'b1110010011010110;
				18'b011000100000011001: oled_data = 16'b1110010011010110;
				18'b011000100010011001: oled_data = 16'b1100001111110010;
				18'b011000100100011001: oled_data = 16'b1101110010010101;
				18'b011000100110011001: oled_data = 16'b1101110011010110;
				18'b011000101000011001: oled_data = 16'b1101110011010101;
				18'b011000101010011001: oled_data = 16'b1101010101110110;
				18'b011000101100011001: oled_data = 16'b1101110111110111;
				18'b011000101110011001: oled_data = 16'b1101010010110100;
				18'b011000110000011001: oled_data = 16'b1101110010110101;
				18'b011000110010011001: oled_data = 16'b1101010010010100;
				18'b011000110100011001: oled_data = 16'b1101110011010110;
				18'b011000110110011001: oled_data = 16'b1101110011010101;
				18'b011000111000011001: oled_data = 16'b1101110011010101;
				18'b011000111010011001: oled_data = 16'b1101110011010101;
				18'b011000111100011001: oled_data = 16'b1101110011010101;
				18'b011000111110011001: oled_data = 16'b1101110011010101;
				18'b011001000000011001: oled_data = 16'b1101110011010101;
				18'b011001000010011001: oled_data = 16'b1101110010110101;
				18'b011001000100011001: oled_data = 16'b1100110000110011;
				18'b011001000110011001: oled_data = 16'b1110010011010110;
				18'b011001001000011001: oled_data = 16'b1110010011010110;
				18'b011001001010011001: oled_data = 16'b1100110000110011;
				18'b011001001100011001: oled_data = 16'b1101010010010100;
				18'b011001001110011001: oled_data = 16'b1101110011010110;
				18'b011001010000011001: oled_data = 16'b1101110011010101;
				18'b011001010010011001: oled_data = 16'b1101110011010101;
				18'b011001010100011001: oled_data = 16'b1101110010110101;
				18'b011001010110011001: oled_data = 16'b1100110000110011;
				18'b011001011000011001: oled_data = 16'b1101110010110101;
				18'b011001011010011001: oled_data = 16'b1110010011010101;
				18'b011001011100011001: oled_data = 16'b1101110011010101;
				18'b011001011110011001: oled_data = 16'b1101110011010101;
				18'b011001100000011001: oled_data = 16'b1110010011010110;
				18'b011001100010011001: oled_data = 16'b1110010011010110;
				18'b011001100100011001: oled_data = 16'b1110010011010110;
				18'b011001100110011001: oled_data = 16'b1101110011010110;
				18'b011001101000011001: oled_data = 16'b1101110011010110;
				18'b011001101010011001: oled_data = 16'b1101110011010110;
				18'b011001101100011001: oled_data = 16'b1101110011010110;
				18'b011001101110011001: oled_data = 16'b1101110011010110;
				18'b011001110000011001: oled_data = 16'b1110010011010110;
				18'b011001110010011001: oled_data = 16'b1101110010110101;
				18'b011001110100011001: oled_data = 16'b1101010001110100;
				18'b011001110110011001: oled_data = 16'b1101110011010101;
				18'b011001111000011001: oled_data = 16'b1101110011010101;
				18'b011001111010011001: oled_data = 16'b1101110011010101;
				18'b011001111100011001: oled_data = 16'b1101110011010101;
				18'b011001111110011001: oled_data = 16'b1101110011010101;
				18'b011010000000011001: oled_data = 16'b1101110011010110;
				18'b011010000010011001: oled_data = 16'b1101010001110100;
				18'b011010000100011001: oled_data = 16'b1110010011110100;
				18'b011010000110011001: oled_data = 16'b1101110001110001;
				18'b011010001000011001: oled_data = 16'b1011101001101010;
				18'b011010001010011001: oled_data = 16'b1011001001001001;
				18'b011010001100011001: oled_data = 16'b1011001001001001;
				18'b011010001110011001: oled_data = 16'b1011001001001001;
				18'b011010010000011001: oled_data = 16'b1011001001001001;
				18'b011010010010011001: oled_data = 16'b1011001001001001;
				18'b011010010100011001: oled_data = 16'b1011001000101001;
				18'b011010010110011001: oled_data = 16'b1010101000001000;
				18'b011010011000011001: oled_data = 16'b1011001001001001;
				18'b011010011010011001: oled_data = 16'b1011001001001001;
				18'b011010011100011001: oled_data = 16'b1011001001001001;
				18'b011010011110011001: oled_data = 16'b1011001000101001;
				18'b011010100000011001: oled_data = 16'b1011001000101001;
				18'b011010100010011001: oled_data = 16'b1011001000101000;
				18'b011010100100011001: oled_data = 16'b1011001000101000;
				18'b011010100110011001: oled_data = 16'b1010101000101000;
				18'b011000011000011010: oled_data = 16'b1110010011110110;
				18'b011000011010011010: oled_data = 16'b1011110001001111;
				18'b011000011100011010: oled_data = 16'b1100110010010010;
				18'b011000011110011010: oled_data = 16'b1101110011010110;
				18'b011000100000011010: oled_data = 16'b1110010011110110;
				18'b011000100010011010: oled_data = 16'b1100001111010010;
				18'b011000100100011010: oled_data = 16'b1101010001110100;
				18'b011000100110011010: oled_data = 16'b1110010011010110;
				18'b011000101000011010: oled_data = 16'b1101110011010101;
				18'b011000101010011010: oled_data = 16'b1101010101110110;
				18'b011000101100011010: oled_data = 16'b1110111010011010;
				18'b011000101110011010: oled_data = 16'b1101010011010101;
				18'b011000110000011010: oled_data = 16'b1101110011010101;
				18'b011000110010011010: oled_data = 16'b1101010001110100;
				18'b011000110100011010: oled_data = 16'b1101110011010110;
				18'b011000110110011010: oled_data = 16'b1110010011010110;
				18'b011000111000011010: oled_data = 16'b1101110011010101;
				18'b011000111010011010: oled_data = 16'b1101110011010101;
				18'b011000111100011010: oled_data = 16'b1101110011010101;
				18'b011000111110011010: oled_data = 16'b1101110011010101;
				18'b011001000000011010: oled_data = 16'b1101110011010101;
				18'b011001000010011010: oled_data = 16'b1101110011010101;
				18'b011001000100011010: oled_data = 16'b1100110000110011;
				18'b011001000110011010: oled_data = 16'b1101110010110101;
				18'b011001001000011010: oled_data = 16'b1101110011010110;
				18'b011001001010011010: oled_data = 16'b1101010010010101;
				18'b011001001100011010: oled_data = 16'b1101010001010100;
				18'b011001001110011010: oled_data = 16'b1101110011010101;
				18'b011001010000011010: oled_data = 16'b1101110011010101;
				18'b011001010010011010: oled_data = 16'b1101110011010101;
				18'b011001010100011010: oled_data = 16'b1101110011010101;
				18'b011001010110011010: oled_data = 16'b1101010010010100;
				18'b011001011000011010: oled_data = 16'b1101010010010100;
				18'b011001011010011010: oled_data = 16'b1101110011010101;
				18'b011001011100011010: oled_data = 16'b1101110011010101;
				18'b011001011110011010: oled_data = 16'b1101110011010101;
				18'b011001100000011010: oled_data = 16'b1101110011010101;
				18'b011001100010011010: oled_data = 16'b1101110011010101;
				18'b011001100100011010: oled_data = 16'b1101110011010101;
				18'b011001100110011010: oled_data = 16'b1101110011010101;
				18'b011001101000011010: oled_data = 16'b1101110011010101;
				18'b011001101010011010: oled_data = 16'b1101110011010101;
				18'b011001101100011010: oled_data = 16'b1101110011010101;
				18'b011001101110011010: oled_data = 16'b1101110011010101;
				18'b011001110000011010: oled_data = 16'b1101110010110101;
				18'b011001110010011010: oled_data = 16'b1101010001010100;
				18'b011001110100011010: oled_data = 16'b1101110010110101;
				18'b011001110110011010: oled_data = 16'b1110010011010110;
				18'b011001111000011010: oled_data = 16'b1101110011010101;
				18'b011001111010011010: oled_data = 16'b1101110011010101;
				18'b011001111100011010: oled_data = 16'b1101110011010110;
				18'b011001111110011010: oled_data = 16'b1101110011010110;
				18'b011010000000011010: oled_data = 16'b1101010010010100;
				18'b011010000010011010: oled_data = 16'b1101110010110100;
				18'b011010000100011010: oled_data = 16'b1110110100010100;
				18'b011010000110011010: oled_data = 16'b1100001101001101;
				18'b011010001000011010: oled_data = 16'b1011001001001001;
				18'b011010001010011010: oled_data = 16'b1011001001001001;
				18'b011010001100011010: oled_data = 16'b1011001001001001;
				18'b011010001110011010: oled_data = 16'b1011001001001001;
				18'b011010010000011010: oled_data = 16'b1011001001001001;
				18'b011010010010011010: oled_data = 16'b1011001001001001;
				18'b011010010100011010: oled_data = 16'b1010101000001000;
				18'b011010010110011010: oled_data = 16'b1011001000101001;
				18'b011010011000011010: oled_data = 16'b1011001001001001;
				18'b011010011010011010: oled_data = 16'b1011001001001001;
				18'b011010011100011010: oled_data = 16'b1011001001001001;
				18'b011010011110011010: oled_data = 16'b1011001000101001;
				18'b011010100000011010: oled_data = 16'b1011001000101001;
				18'b011010100010011010: oled_data = 16'b1011001000101000;
				18'b011010100100011010: oled_data = 16'b1011001000101000;
				18'b011010100110011010: oled_data = 16'b1010101000101000;
				18'b011000011000011011: oled_data = 16'b1101110011010110;
				18'b011000011010011011: oled_data = 16'b1011010001001100;
				18'b011000011100011011: oled_data = 16'b1100110010010001;
				18'b011000011110011011: oled_data = 16'b1101110011010110;
				18'b011000100000011011: oled_data = 16'b1110010011010110;
				18'b011000100010011011: oled_data = 16'b1100010000010010;
				18'b011000100100011011: oled_data = 16'b1101010001010100;
				18'b011000100110011011: oled_data = 16'b1110010011110110;
				18'b011000101000011011: oled_data = 16'b1101110010110101;
				18'b011000101010011011: oled_data = 16'b1101110110110111;
				18'b011000101100011011: oled_data = 16'b1110111011011010;
				18'b011000101110011011: oled_data = 16'b1101010101010110;
				18'b011000110000011011: oled_data = 16'b1101110010110101;
				18'b011000110010011011: oled_data = 16'b1101010001110100;
				18'b011000110100011011: oled_data = 16'b1101110011010101;
				18'b011000110110011011: oled_data = 16'b1110010011010110;
				18'b011000111000011011: oled_data = 16'b1101110011010101;
				18'b011000111010011011: oled_data = 16'b1101110011010101;
				18'b011000111100011011: oled_data = 16'b1110010011010110;
				18'b011000111110011011: oled_data = 16'b1110010011010110;
				18'b011001000000011011: oled_data = 16'b1101110011010101;
				18'b011001000010011011: oled_data = 16'b1101110011010110;
				18'b011001000100011011: oled_data = 16'b1100110001110100;
				18'b011001000110011011: oled_data = 16'b1101010010010100;
				18'b011001001000011011: oled_data = 16'b1101110011010110;
				18'b011001001010011011: oled_data = 16'b1101110011010101;
				18'b011001001100011011: oled_data = 16'b1101010001110100;
				18'b011001001110011011: oled_data = 16'b1101010010110101;
				18'b011001010000011011: oled_data = 16'b1101110011010101;
				18'b011001010010011011: oled_data = 16'b1101110011010101;
				18'b011001010100011011: oled_data = 16'b1101110011010101;
				18'b011001010110011011: oled_data = 16'b1101110010110101;
				18'b011001011000011011: oled_data = 16'b1101010100010101;
				18'b011001011010011011: oled_data = 16'b1101010011010101;
				18'b011001011100011011: oled_data = 16'b1110010011010101;
				18'b011001011110011011: oled_data = 16'b1101110011010101;
				18'b011001100000011011: oled_data = 16'b1101110011010101;
				18'b011001100010011011: oled_data = 16'b1101110011010110;
				18'b011001100100011011: oled_data = 16'b1101110011010110;
				18'b011001100110011011: oled_data = 16'b1110010011010110;
				18'b011001101000011011: oled_data = 16'b1110010011110110;
				18'b011001101010011011: oled_data = 16'b1110010011110110;
				18'b011001101100011011: oled_data = 16'b1101110011010101;
				18'b011001101110011011: oled_data = 16'b1101010011010101;
				18'b011001110000011011: oled_data = 16'b1100010100010100;
				18'b011001110010011011: oled_data = 16'b1100110011110101;
				18'b011001110100011011: oled_data = 16'b1101110011010101;
				18'b011001110110011011: oled_data = 16'b1101110011010101;
				18'b011001111000011011: oled_data = 16'b1101110011010101;
				18'b011001111010011011: oled_data = 16'b1101110010110101;
				18'b011001111100011011: oled_data = 16'b1101010001110100;
				18'b011001111110011011: oled_data = 16'b1101010010110101;
				18'b011010000000011011: oled_data = 16'b1100110001010010;
				18'b011010000010011011: oled_data = 16'b1110010011110100;
				18'b011010000100011011: oled_data = 16'b1101110001110001;
				18'b011010000110011011: oled_data = 16'b1011001001101001;
				18'b011010001000011011: oled_data = 16'b1011101001001001;
				18'b011010001010011011: oled_data = 16'b1100001011001100;
				18'b011010001100011011: oled_data = 16'b1011101001101010;
				18'b011010001110011011: oled_data = 16'b1011001001001001;
				18'b011010010000011011: oled_data = 16'b1011101001001001;
				18'b011010010010011011: oled_data = 16'b1011001000101000;
				18'b011010010100011011: oled_data = 16'b1010101000101001;
				18'b011010010110011011: oled_data = 16'b1011001001001001;
				18'b011010011000011011: oled_data = 16'b1011001001001001;
				18'b011010011010011011: oled_data = 16'b1011001000101001;
				18'b011010011100011011: oled_data = 16'b1011001000101001;
				18'b011010011110011011: oled_data = 16'b1011001000101001;
				18'b011010100000011011: oled_data = 16'b1011001000101001;
				18'b011010100010011011: oled_data = 16'b1011001000101000;
				18'b011010100100011011: oled_data = 16'b1011001000101000;
				18'b011010100110011011: oled_data = 16'b1010101000101000;
				18'b011000011000011100: oled_data = 16'b1101110010110110;
				18'b011000011010011100: oled_data = 16'b1011010000101011;
				18'b011000011100011100: oled_data = 16'b1100110001110000;
				18'b011000011110011100: oled_data = 16'b1110010011010110;
				18'b011000100000011100: oled_data = 16'b1110010011010110;
				18'b011000100010011100: oled_data = 16'b1100010000010010;
				18'b011000100100011100: oled_data = 16'b1100110000010011;
				18'b011000100110011100: oled_data = 16'b1110010011110110;
				18'b011000101000011100: oled_data = 16'b1101110010110101;
				18'b011000101010011100: oled_data = 16'b1101010110110111;
				18'b011000101100011100: oled_data = 16'b1110011010111010;
				18'b011000101110011100: oled_data = 16'b1101111000111000;
				18'b011000110000011100: oled_data = 16'b1101010011010101;
				18'b011000110010011100: oled_data = 16'b1101010010010100;
				18'b011000110100011100: oled_data = 16'b1101110010010101;
				18'b011000110110011100: oled_data = 16'b1101110011010110;
				18'b011000111000011100: oled_data = 16'b1101110011010101;
				18'b011000111010011100: oled_data = 16'b1101110011010101;
				18'b011000111100011100: oled_data = 16'b1110010011010110;
				18'b011000111110011100: oled_data = 16'b1110010011010110;
				18'b011001000000011100: oled_data = 16'b1101110011010101;
				18'b011001000010011100: oled_data = 16'b1101110011010110;
				18'b011001000100011100: oled_data = 16'b1101010011010101;
				18'b011001000110011100: oled_data = 16'b1100110011010100;
				18'b011001001000011100: oled_data = 16'b1101010011010101;
				18'b011001001010011100: oled_data = 16'b1110010011010101;
				18'b011001001100011100: oled_data = 16'b1101010010110100;
				18'b011001001110011100: oled_data = 16'b1100110010110100;
				18'b011001010000011100: oled_data = 16'b1101110011010101;
				18'b011001010010011100: oled_data = 16'b1101110011010110;
				18'b011001010100011100: oled_data = 16'b1101110011010101;
				18'b011001010110011100: oled_data = 16'b1101110010110101;
				18'b011001011000011100: oled_data = 16'b1101110111011000;
				18'b011001011010011100: oled_data = 16'b1101010110110111;
				18'b011001011100011100: oled_data = 16'b1101010010110100;
				18'b011001011110011100: oled_data = 16'b1101110011010110;
				18'b011001100000011100: oled_data = 16'b1101110011010101;
				18'b011001100010011100: oled_data = 16'b1101010001010100;
				18'b011001100100011100: oled_data = 16'b1100110000110011;
				18'b011001100110011100: oled_data = 16'b1100110000110011;
				18'b011001101000011100: oled_data = 16'b1100110000110011;
				18'b011001101010011100: oled_data = 16'b1100110000010011;
				18'b011001101100011100: oled_data = 16'b1100001111110010;
				18'b011001101110011100: oled_data = 16'b1101010011010101;
				18'b011001110000011100: oled_data = 16'b1110111011111011;
				18'b011001110010011100: oled_data = 16'b1110111011111011;
				18'b011001110100011100: oled_data = 16'b1101010110010110;
				18'b011001110110011100: oled_data = 16'b1101010010110101;
				18'b011001111000011100: oled_data = 16'b1110010011010110;
				18'b011001111010011100: oled_data = 16'b1110010011110110;
				18'b011001111100011100: oled_data = 16'b1101010010010100;
				18'b011001111110011100: oled_data = 16'b1100010000110011;
				18'b011010000000011100: oled_data = 16'b1100110001010010;
				18'b011010000010011100: oled_data = 16'b1110110100010100;
				18'b011010000100011100: oled_data = 16'b1100101101101110;
				18'b011010000110011100: oled_data = 16'b1011001000101001;
				18'b011010001000011100: oled_data = 16'b1011101010001010;
				18'b011010001010011100: oled_data = 16'b1101001110001110;
				18'b011010001100011100: oled_data = 16'b1011001001001010;
				18'b011010001110011100: oled_data = 16'b1011001001001001;
				18'b011010010000011100: oled_data = 16'b1011001001001001;
				18'b011010010010011100: oled_data = 16'b1010101000001000;
				18'b011010010100011100: oled_data = 16'b1011101001001001;
				18'b011010010110011100: oled_data = 16'b1011001001001001;
				18'b011010011000011100: oled_data = 16'b1010000111101000;
				18'b011010011010011100: oled_data = 16'b1010000111000111;
				18'b011010011100011100: oled_data = 16'b1011001001001001;
				18'b011010011110011100: oled_data = 16'b1011001000101001;
				18'b011010100000011100: oled_data = 16'b1011001000101001;
				18'b011010100010011100: oled_data = 16'b1011001000101000;
				18'b011010100100011100: oled_data = 16'b1011001000101000;
				18'b011010100110011100: oled_data = 16'b1010101000101000;
				18'b011000011000011101: oled_data = 16'b1101110010110101;
				18'b011000011010011101: oled_data = 16'b1010110000101010;
				18'b011000011100011101: oled_data = 16'b1100010010001110;
				18'b011000011110011101: oled_data = 16'b1110010011010110;
				18'b011000100000011101: oled_data = 16'b1110010011010110;
				18'b011000100010011101: oled_data = 16'b1100110000110011;
				18'b011000100100011101: oled_data = 16'b1011101111010001;
				18'b011000100110011101: oled_data = 16'b1110010011110110;
				18'b011000101000011101: oled_data = 16'b1101110010110101;
				18'b011000101010011101: oled_data = 16'b1101010110010110;
				18'b011000101100011101: oled_data = 16'b1110111100011011;
				18'b011000101110011101: oled_data = 16'b1101111001011001;
				18'b011000110000011101: oled_data = 16'b1100110100010101;
				18'b011000110010011101: oled_data = 16'b1101110010110101;
				18'b011000110100011101: oled_data = 16'b1101010001110100;
				18'b011000110110011101: oled_data = 16'b1101110011010110;
				18'b011000111000011101: oled_data = 16'b1101110011010101;
				18'b011000111010011101: oled_data = 16'b1101110011010101;
				18'b011000111100011101: oled_data = 16'b1101110011010110;
				18'b011000111110011101: oled_data = 16'b1101110011010110;
				18'b011001000000011101: oled_data = 16'b1101110011010101;
				18'b011001000010011101: oled_data = 16'b1101110011010101;
				18'b011001000100011101: oled_data = 16'b1101110011010101;
				18'b011001000110011101: oled_data = 16'b1101010110010110;
				18'b011001001000011101: oled_data = 16'b1101010011010101;
				18'b011001001010011101: oled_data = 16'b1101110011010101;
				18'b011001001100011101: oled_data = 16'b1101110011010101;
				18'b011001001110011101: oled_data = 16'b1101010100110110;
				18'b011001010000011101: oled_data = 16'b1101010010110101;
				18'b011001010010011101: oled_data = 16'b1101110010010101;
				18'b011001010100011101: oled_data = 16'b1101110010110101;
				18'b011001010110011101: oled_data = 16'b1101110011010101;
				18'b011001011000011101: oled_data = 16'b1101010101010110;
				18'b011001011010011101: oled_data = 16'b1110111011111011;
				18'b011001011100011101: oled_data = 16'b1101110101110110;
				18'b011001011110011101: oled_data = 16'b1101110010110101;
				18'b011001100000011101: oled_data = 16'b1101110011010110;
				18'b011001100010011101: oled_data = 16'b1101010010010100;
				18'b011001100100011101: oled_data = 16'b1011001110010000;
				18'b011001100110011101: oled_data = 16'b1011001101110000;
				18'b011001101000011101: oled_data = 16'b1011101110110001;
				18'b011001101010011101: oled_data = 16'b1100110001010011;
				18'b011001101100011101: oled_data = 16'b1101110010110101;
				18'b011001101110011101: oled_data = 16'b1101110011010101;
				18'b011001110000011101: oled_data = 16'b1101010110010110;
				18'b011001110010011101: oled_data = 16'b1101111001111000;
				18'b011001110100011101: oled_data = 16'b1110011010111010;
				18'b011001110110011101: oled_data = 16'b1011110001010011;
				18'b011001111000011101: oled_data = 16'b1100101111110011;
				18'b011001111010011101: oled_data = 16'b1101010001010100;
				18'b011001111100011101: oled_data = 16'b1100010000110011;
				18'b011001111110011101: oled_data = 16'b1011001110110000;
				18'b011010000000011101: oled_data = 16'b1101110011010011;
				18'b011010000010011101: oled_data = 16'b1110010011010011;
				18'b011010000100011101: oled_data = 16'b1011101010101011;
				18'b011010000110011101: oled_data = 16'b1011001000101001;
				18'b011010001000011101: oled_data = 16'b1100001011101011;
				18'b011010001010011101: oled_data = 16'b1100001100001100;
				18'b011010001100011101: oled_data = 16'b1011001000101001;
				18'b011010001110011101: oled_data = 16'b1011001001001001;
				18'b011010010000011101: oled_data = 16'b1010101000101000;
				18'b011010010010011101: oled_data = 16'b1011001001001001;
				18'b011010010100011101: oled_data = 16'b1011101001001010;
				18'b011010010110011101: oled_data = 16'b1010001000001000;
				18'b011010011000011101: oled_data = 16'b1001000101100110;
				18'b011010011010011101: oled_data = 16'b1010101000001000;
				18'b011010011100011101: oled_data = 16'b1011001000101001;
				18'b011010011110011101: oled_data = 16'b1011001000101001;
				18'b011010100000011101: oled_data = 16'b1011001000101001;
				18'b011010100010011101: oled_data = 16'b1011001000101000;
				18'b011010100100011101: oled_data = 16'b1011001000101000;
				18'b011010100110011101: oled_data = 16'b1010101000101000;
				18'b011000011000011110: oled_data = 16'b1101110010110101;
				18'b011000011010011110: oled_data = 16'b1011010001001001;
				18'b011000011100011110: oled_data = 16'b1011110001101100;
				18'b011000011110011110: oled_data = 16'b1101110011010110;
				18'b011000100000011110: oled_data = 16'b1101110011010110;
				18'b011000100010011110: oled_data = 16'b1101010001110100;
				18'b011000100100011110: oled_data = 16'b1011101110110001;
				18'b011000100110011110: oled_data = 16'b1101110011010110;
				18'b011000101000011110: oled_data = 16'b1101110010110101;
				18'b011000101010011110: oled_data = 16'b1101010101010110;
				18'b011000101100011110: oled_data = 16'b1110111100011011;
				18'b011000101110011110: oled_data = 16'b1110111011011010;
				18'b011000110000011110: oled_data = 16'b1101010101010110;
				18'b011000110010011110: oled_data = 16'b1101110010110101;
				18'b011000110100011110: oled_data = 16'b1101010001110100;
				18'b011000110110011110: oled_data = 16'b1101110011010101;
				18'b011000111000011110: oled_data = 16'b1101110011010101;
				18'b011000111010011110: oled_data = 16'b1101110011010101;
				18'b011000111100011110: oled_data = 16'b1101110011010101;
				18'b011000111110011110: oled_data = 16'b1101110011010101;
				18'b011001000000011110: oled_data = 16'b1101110011010101;
				18'b011001000010011110: oled_data = 16'b1101110011010101;
				18'b011001000100011110: oled_data = 16'b1101110010110101;
				18'b011001000110011110: oled_data = 16'b1101110111111000;
				18'b011001001000011110: oled_data = 16'b1101110110110111;
				18'b011001001010011110: oled_data = 16'b1101110011010101;
				18'b011001001100011110: oled_data = 16'b1101110011010101;
				18'b011001001110011110: oled_data = 16'b1101110111011000;
				18'b011001010000011110: oled_data = 16'b1100010011010100;
				18'b011001010010011110: oled_data = 16'b1101010001110100;
				18'b011001010100011110: oled_data = 16'b1101110011010110;
				18'b011001010110011110: oled_data = 16'b1101110011010101;
				18'b011001011000011110: oled_data = 16'b1101010011110101;
				18'b011001011010011110: oled_data = 16'b1110011010011010;
				18'b011001011100011110: oled_data = 16'b1110011011111011;
				18'b011001011110011110: oled_data = 16'b1101010101010110;
				18'b011001100000011110: oled_data = 16'b1101110011010101;
				18'b011001100010011110: oled_data = 16'b1101110011110110;
				18'b011001100100011110: oled_data = 16'b1101010001010100;
				18'b011001100110011110: oled_data = 16'b1100110001010011;
				18'b011001101000011110: oled_data = 16'b1101110011010101;
				18'b011001101010011110: oled_data = 16'b1101110011010110;
				18'b011001101100011110: oled_data = 16'b1101110011010101;
				18'b011001101110011110: oled_data = 16'b1110010011010110;
				18'b011001110000011110: oled_data = 16'b1100110010110100;
				18'b011001110010011110: oled_data = 16'b1100110110110101;
				18'b011001110100011110: oled_data = 16'b1110111011111010;
				18'b011001110110011110: oled_data = 16'b1100110100110101;
				18'b011001111000011110: oled_data = 16'b1011001101110000;
				18'b011001111010011110: oled_data = 16'b1011001110010001;
				18'b011001111100011110: oled_data = 16'b1011001101110000;
				18'b011001111110011110: oled_data = 16'b1100001111110001;
				18'b011010000000011110: oled_data = 16'b1110110100010100;
				18'b011010000010011110: oled_data = 16'b1101001111110000;
				18'b011010000100011110: oled_data = 16'b1011001000101001;
				18'b011010000110011110: oled_data = 16'b1011001001001001;
				18'b011010001000011110: oled_data = 16'b1100001100001100;
				18'b011010001010011110: oled_data = 16'b1011101010001010;
				18'b011010001100011110: oled_data = 16'b1011001001001001;
				18'b011010001110011110: oled_data = 16'b1011001001001001;
				18'b011010010000011110: oled_data = 16'b1010101000101000;
				18'b011010010010011110: oled_data = 16'b1011001001001001;
				18'b011010010100011110: oled_data = 16'b1010101000101000;
				18'b011010010110011110: oled_data = 16'b1000100101100110;
				18'b011010011000011110: oled_data = 16'b1001100110100111;
				18'b011010011010011110: oled_data = 16'b1011101010001011;
				18'b011010011100011110: oled_data = 16'b1011101010101010;
				18'b011010011110011110: oled_data = 16'b1011001000101000;
				18'b011010100000011110: oled_data = 16'b1011001000101001;
				18'b011010100010011110: oled_data = 16'b1011001000101000;
				18'b011010100100011110: oled_data = 16'b1011001000101000;
				18'b011010100110011110: oled_data = 16'b1010101000101000;
				18'b011000011000011111: oled_data = 16'b1101010010110101;
				18'b011000011010011111: oled_data = 16'b1011010001101001;
				18'b011000011100011111: oled_data = 16'b1011010001001011;
				18'b011000011110011111: oled_data = 16'b1101110010110101;
				18'b011000100000011111: oled_data = 16'b1101110011010110;
				18'b011000100010011111: oled_data = 16'b1101010010010100;
				18'b011000100100011111: oled_data = 16'b1011001101110000;
				18'b011000100110011111: oled_data = 16'b1101110010110101;
				18'b011000101000011111: oled_data = 16'b1101110010110101;
				18'b011000101010011111: oled_data = 16'b1101010101010110;
				18'b011000101100011111: oled_data = 16'b1110111100011011;
				18'b011000101110011111: oled_data = 16'b1110111100011011;
				18'b011000110000011111: oled_data = 16'b1101111000111001;
				18'b011000110010011111: oled_data = 16'b1100110010010100;
				18'b011000110100011111: oled_data = 16'b1101110010110101;
				18'b011000110110011111: oled_data = 16'b1101110010010101;
				18'b011000111000011111: oled_data = 16'b1101110011010110;
				18'b011000111010011111: oled_data = 16'b1101110011010101;
				18'b011000111100011111: oled_data = 16'b1101110011010101;
				18'b011000111110011111: oled_data = 16'b1101110011010101;
				18'b011001000000011111: oled_data = 16'b1101110011010101;
				18'b011001000010011111: oled_data = 16'b1101110011010101;
				18'b011001000100011111: oled_data = 16'b1101110011010101;
				18'b011001000110011111: oled_data = 16'b1101110101110111;
				18'b011001001000011111: oled_data = 16'b1101111010011001;
				18'b011001001010011111: oled_data = 16'b1100110010110100;
				18'b011001001100011111: oled_data = 16'b1101010001110100;
				18'b011001001110011111: oled_data = 16'b1101010101110110;
				18'b011001010000011111: oled_data = 16'b1110011010011010;
				18'b011001010010011111: oled_data = 16'b1101010011110101;
				18'b011001010100011111: oled_data = 16'b1101110011010101;
				18'b011001010110011111: oled_data = 16'b1101110011010101;
				18'b011001011000011111: oled_data = 16'b1101110010110101;
				18'b011001011010011111: oled_data = 16'b1101110111110111;
				18'b011001011100011111: oled_data = 16'b1110111100111011;
				18'b011001011110011111: oled_data = 16'b1110111011011010;
				18'b011001100000011111: oled_data = 16'b1100010010110100;
				18'b011001100010011111: oled_data = 16'b1101110010110101;
				18'b011001100100011111: oled_data = 16'b1101110011010101;
				18'b011001100110011111: oled_data = 16'b1101010010010100;
				18'b011001101000011111: oled_data = 16'b1101010010010100;
				18'b011001101010011111: oled_data = 16'b1101110011010101;
				18'b011001101100011111: oled_data = 16'b1101110011010101;
				18'b011001101110011111: oled_data = 16'b1101110011010101;
				18'b011001110000011111: oled_data = 16'b1101110011010101;
				18'b011001110010011111: oled_data = 16'b1101010100110101;
				18'b011001110100011111: oled_data = 16'b1110111010111010;
				18'b011001110110011111: oled_data = 16'b1101010111011000;
				18'b011001111000011111: oled_data = 16'b1011001110010001;
				18'b011001111010011111: oled_data = 16'b1011001110010001;
				18'b011001111100011111: oled_data = 16'b1010101101101111;
				18'b011001111110011111: oled_data = 16'b1101010010010010;
				18'b011010000000011111: oled_data = 16'b1110110100010100;
				18'b011010000010011111: oled_data = 16'b1011101100001101;
				18'b011010000100011111: oled_data = 16'b1011001000101001;
				18'b011010000110011111: oled_data = 16'b1011101001001001;
				18'b011010001000011111: oled_data = 16'b1011101010001010;
				18'b011010001010011111: oled_data = 16'b1011001001001001;
				18'b011010001100011111: oled_data = 16'b1011001001001001;
				18'b011010001110011111: oled_data = 16'b1010101000101000;
				18'b011010010000011111: oled_data = 16'b1011001001001001;
				18'b011010010010011111: oled_data = 16'b1011001000101001;
				18'b011010010100011111: oled_data = 16'b1001000110000111;
				18'b011010010110011111: oled_data = 16'b1001000101100110;
				18'b011010011000011111: oled_data = 16'b1011001001001001;
				18'b011010011010011111: oled_data = 16'b1101001111101111;
				18'b011010011100011111: oled_data = 16'b1011101010001010;
				18'b011010011110011111: oled_data = 16'b1011001000101000;
				18'b011010100000011111: oled_data = 16'b1011001000101001;
				18'b011010100010011111: oled_data = 16'b1011001000101000;
				18'b011010100100011111: oled_data = 16'b1011001000101000;
				18'b011010100110011111: oled_data = 16'b1010101000001000;
				18'b011000011000100000: oled_data = 16'b1101010001110101;
				18'b011000011010100000: oled_data = 16'b1011010001101001;
				18'b011000011100100000: oled_data = 16'b1011110001101100;
				18'b011000011110100000: oled_data = 16'b1101010010010101;
				18'b011000100000100000: oled_data = 16'b1101110011010110;
				18'b011000100010100000: oled_data = 16'b1101110010110101;
				18'b011000100100100000: oled_data = 16'b1011001110010001;
				18'b011000100110100000: oled_data = 16'b1101010001110100;
				18'b011000101000100000: oled_data = 16'b1101110011010110;
				18'b011000101010100000: oled_data = 16'b1010110000010001;
				18'b011000101100100000: oled_data = 16'b1101011001011000;
				18'b011000101110100000: oled_data = 16'b1110111100111011;
				18'b011000110000100000: oled_data = 16'b1110111011111011;
				18'b011000110010100000: oled_data = 16'b1100110101010110;
				18'b011000110100100000: oled_data = 16'b1101010010010100;
				18'b011000110110100000: oled_data = 16'b1101010001010100;
				18'b011000111000100000: oled_data = 16'b1101110011010101;
				18'b011000111010100000: oled_data = 16'b1101110011010101;
				18'b011000111100100000: oled_data = 16'b1101110011010101;
				18'b011000111110100000: oled_data = 16'b1101110011010101;
				18'b011001000000100000: oled_data = 16'b1101110010110101;
				18'b011001000010100000: oled_data = 16'b1101110010110101;
				18'b011001000100100000: oled_data = 16'b1101110010110101;
				18'b011001000110100000: oled_data = 16'b1100110011010100;
				18'b011001001000100000: oled_data = 16'b1101011010011000;
				18'b011001001010100000: oled_data = 16'b1100110100010101;
				18'b011001001100100000: oled_data = 16'b1101110010110101;
				18'b011001001110100000: oled_data = 16'b1101010101010110;
				18'b011001010000100000: oled_data = 16'b1110111100011011;
				18'b011001010010100000: oled_data = 16'b1110011001011001;
				18'b011001010100100000: oled_data = 16'b1101010011110101;
				18'b011001010110100000: oled_data = 16'b1110010011110110;
				18'b011001011000100000: oled_data = 16'b1101110010110100;
				18'b011001011010100000: oled_data = 16'b1100010011010011;
				18'b011001011100100000: oled_data = 16'b1110111100011010;
				18'b011001011110100000: oled_data = 16'b1110111100111011;
				18'b011001100000100000: oled_data = 16'b1100110110010110;
				18'b011001100010100000: oled_data = 16'b1011101111010001;
				18'b011001100100100000: oled_data = 16'b1101110010110101;
				18'b011001100110100000: oled_data = 16'b1110010011110110;
				18'b011001101000100000: oled_data = 16'b1101010010010100;
				18'b011001101010100000: oled_data = 16'b1101010001110100;
				18'b011001101100100000: oled_data = 16'b1101110011010101;
				18'b011001101110100000: oled_data = 16'b1101110011110110;
				18'b011001110000100000: oled_data = 16'b1101110011010101;
				18'b011001110010100000: oled_data = 16'b1101110011010101;
				18'b011001110100100000: oled_data = 16'b1101010110010111;
				18'b011001110110100000: oled_data = 16'b1101010111111000;
				18'b011001111000100000: oled_data = 16'b1011001110010001;
				18'b011001111010100000: oled_data = 16'b1011001101110000;
				18'b011001111100100000: oled_data = 16'b1011001110010000;
				18'b011001111110100000: oled_data = 16'b1101110011110011;
				18'b011010000000100000: oled_data = 16'b1110010011110011;
				18'b011010000010100000: oled_data = 16'b1011001001101010;
				18'b011010000100100000: oled_data = 16'b1011001000101001;
				18'b011010000110100000: oled_data = 16'b1011001001001001;
				18'b011010001000100000: oled_data = 16'b1011001001001001;
				18'b011010001010100000: oled_data = 16'b1011001001001001;
				18'b011010001100100000: oled_data = 16'b1011001001001001;
				18'b011010001110100000: oled_data = 16'b1010101000101001;
				18'b011010010000100000: oled_data = 16'b1011001001001001;
				18'b011010010010100000: oled_data = 16'b1001100110100111;
				18'b011010010100100000: oled_data = 16'b1000100101000110;
				18'b011010010110100000: oled_data = 16'b1010000111001000;
				18'b011010011000100000: oled_data = 16'b1100101100101101;
				18'b011010011010100000: oled_data = 16'b1100001100001100;
				18'b011010011100100000: oled_data = 16'b1011001000101000;
				18'b011010011110100000: oled_data = 16'b1011001000101001;
				18'b011010100000100000: oled_data = 16'b1011001000101001;
				18'b011010100010100000: oled_data = 16'b1011001000101000;
				18'b011010100100100000: oled_data = 16'b1011001000101000;
				18'b011010100110100000: oled_data = 16'b1011001000001000;
				18'b011000011000100001: oled_data = 16'b1100110010110010;
				18'b011000011010100001: oled_data = 16'b1011010010001011;
				18'b011000011100100001: oled_data = 16'b1100110010110001;
				18'b011000011110100001: oled_data = 16'b1101010001110100;
				18'b011000100000100001: oled_data = 16'b1101110011010101;
				18'b011000100010100001: oled_data = 16'b1101110011010101;
				18'b011000100100100001: oled_data = 16'b1011101110010001;
				18'b011000100110100001: oled_data = 16'b1100010000010010;
				18'b011000101000100001: oled_data = 16'b1110010100010110;
				18'b011000101010100001: oled_data = 16'b1000001011001100;
				18'b011000101100100001: oled_data = 16'b0101001001001000;
				18'b011000101110100001: oled_data = 16'b1101011000110111;
				18'b011000110000100001: oled_data = 16'b1110111100111011;
				18'b011000110010100001: oled_data = 16'b1101111010011001;
				18'b011000110100100001: oled_data = 16'b1100110011010100;
				18'b011000110110100001: oled_data = 16'b1101010010010100;
				18'b011000111000100001: oled_data = 16'b1101110010110101;
				18'b011000111010100001: oled_data = 16'b1101110011010101;
				18'b011000111100100001: oled_data = 16'b1101110011010110;
				18'b011000111110100001: oled_data = 16'b1101010010010100;
				18'b011001000000100001: oled_data = 16'b1100110001010011;
				18'b011001000010100001: oled_data = 16'b1101010001010100;
				18'b011001000100100001: oled_data = 16'b1101010010010100;
				18'b011001000110100001: oled_data = 16'b1100110011010100;
				18'b011001001000100001: oled_data = 16'b1110011011111010;
				18'b011001001010100001: oled_data = 16'b1101111000111001;
				18'b011001001100100001: oled_data = 16'b1101010011010101;
				18'b011001001110100001: oled_data = 16'b1101010011110101;
				18'b011001010000100001: oled_data = 16'b1110011010111010;
				18'b011001010010100001: oled_data = 16'b1111011101011011;
				18'b011001010100100001: oled_data = 16'b1101111000111000;
				18'b011001010110100001: oled_data = 16'b1001101110101111;
				18'b011001011000100001: oled_data = 16'b0111001000101010;
				18'b011001011010100001: oled_data = 16'b1000101100001101;
				18'b011001011100100001: oled_data = 16'b1110011010011001;
				18'b011001011110100001: oled_data = 16'b1110111100111011;
				18'b011001100000100001: oled_data = 16'b1110011010011010;
				18'b011001100010100001: oled_data = 16'b1010101110110000;
				18'b011001100100100001: oled_data = 16'b1011001110010001;
				18'b011001100110100001: oled_data = 16'b1100001111110010;
				18'b011001101000100001: oled_data = 16'b1101010001110100;
				18'b011001101010100001: oled_data = 16'b1101010001010100;
				18'b011001101100100001: oled_data = 16'b1100110001010011;
				18'b011001101110100001: oled_data = 16'b1101010001110100;
				18'b011001110000100001: oled_data = 16'b1101010010010101;
				18'b011001110010100001: oled_data = 16'b1101110011010101;
				18'b011001110100100001: oled_data = 16'b1101010011010101;
				18'b011001110110100001: oled_data = 16'b1100010011110101;
				18'b011001111000100001: oled_data = 16'b1010101101110000;
				18'b011001111010100001: oled_data = 16'b1010101101010000;
				18'b011001111100100001: oled_data = 16'b1011101111010001;
				18'b011001111110100001: oled_data = 16'b1110010100010100;
				18'b011010000000100001: oled_data = 16'b1101110001110001;
				18'b011010000010100001: oled_data = 16'b1011001000101001;
				18'b011010000100100001: oled_data = 16'b1011101001001001;
				18'b011010000110100001: oled_data = 16'b1011001001001001;
				18'b011010001000100001: oled_data = 16'b1011001001001001;
				18'b011010001010100001: oled_data = 16'b1011001001001001;
				18'b011010001100100001: oled_data = 16'b1010101000101000;
				18'b011010001110100001: oled_data = 16'b1011001001001001;
				18'b011010010000100001: oled_data = 16'b1010000111101000;
				18'b011010010010100001: oled_data = 16'b1000100101000110;
				18'b011010010100100001: oled_data = 16'b1001100110000111;
				18'b011010010110100001: oled_data = 16'b1011001000101001;
				18'b011010011000100001: oled_data = 16'b1011101010001010;
				18'b011010011010100001: oled_data = 16'b1011001001001001;
				18'b011010011100100001: oled_data = 16'b1011001000101001;
				18'b011010011110100001: oled_data = 16'b1011001000101001;
				18'b011010100000100001: oled_data = 16'b1011001000101001;
				18'b011010100010100001: oled_data = 16'b1011001000101000;
				18'b011010100100100001: oled_data = 16'b1011001000101000;
				18'b011010100110100001: oled_data = 16'b1010101000001000;
				18'b011000011000100010: oled_data = 16'b1010010001001111;
				18'b011000011010100010: oled_data = 16'b1010110000101101;
				18'b011000011100100010: oled_data = 16'b1101110010110100;
				18'b011000011110100010: oled_data = 16'b1101010001010100;
				18'b011000100000100010: oled_data = 16'b1101010010010100;
				18'b011000100010100010: oled_data = 16'b1101110011010110;
				18'b011000100100100010: oled_data = 16'b1100001111010010;
				18'b011000100110100010: oled_data = 16'b1011001101110000;
				18'b011000101000100010: oled_data = 16'b1101110011010110;
				18'b011000101010100010: oled_data = 16'b1010101111110001;
				18'b011000101100100010: oled_data = 16'b0011100101000100;
				18'b011000101110100010: oled_data = 16'b0101001000100111;
				18'b011000110000100010: oled_data = 16'b1100111000010111;
				18'b011000110010100010: oled_data = 16'b1110111100111011;
				18'b011000110100100010: oled_data = 16'b1101010110110110;
				18'b011000110110100010: oled_data = 16'b1101110010110101;
				18'b011000111000100010: oled_data = 16'b1101010010010100;
				18'b011000111010100010: oled_data = 16'b1101110011010101;
				18'b011000111100100010: oled_data = 16'b1101110011010110;
				18'b011000111110100010: oled_data = 16'b1101110011010110;
				18'b011001000000100010: oled_data = 16'b1110010011010110;
				18'b011001000010100010: oled_data = 16'b1110010011010110;
				18'b011001000100100010: oled_data = 16'b1110010011010110;
				18'b011001000110100010: oled_data = 16'b1101010011010100;
				18'b011001001000100010: oled_data = 16'b1110011010011001;
				18'b011001001010100010: oled_data = 16'b1110011011111011;
				18'b011001001100100010: oled_data = 16'b1101010100010110;
				18'b011001001110100010: oled_data = 16'b1101110010110101;
				18'b011001010000100010: oled_data = 16'b1110011001111001;
				18'b011001010010100010: oled_data = 16'b1100010111010110;
				18'b011001010100100010: oled_data = 16'b0110001011001011;
				18'b011001010110100010: oled_data = 16'b0011000100100100;
				18'b011001011000100010: oled_data = 16'b0101001000001000;
				18'b011001011010100010: oled_data = 16'b1010001110110000;
				18'b011001011100100010: oled_data = 16'b1101110111010111;
				18'b011001011110100010: oled_data = 16'b1110111100011011;
				18'b011001100000100010: oled_data = 16'b1110111100111011;
				18'b011001100010100010: oled_data = 16'b1100110100010101;
				18'b011001100100100010: oled_data = 16'b1011001101010000;
				18'b011001100110100010: oled_data = 16'b1011001101110001;
				18'b011001101000100010: oled_data = 16'b1011001101110001;
				18'b011001101010100010: oled_data = 16'b1011101110110001;
				18'b011001101100100010: oled_data = 16'b1100010000010011;
				18'b011001101110100010: oled_data = 16'b1100110000110011;
				18'b011001110000100010: oled_data = 16'b1100110001010100;
				18'b011001110010100010: oled_data = 16'b1101110011010101;
				18'b011001110100100010: oled_data = 16'b1101110011010101;
				18'b011001110110100010: oled_data = 16'b1101110010110101;
				18'b011001111000100010: oled_data = 16'b1100010000110011;
				18'b011001111010100010: oled_data = 16'b1011101111010001;
				18'b011001111100100010: oled_data = 16'b1011101111010001;
				18'b011001111110100010: oled_data = 16'b1110110100110100;
				18'b011010000000100010: oled_data = 16'b1100101111001111;
				18'b011010000010100010: oled_data = 16'b1011001000001000;
				18'b011010000100100010: oled_data = 16'b1011101001001001;
				18'b011010000110100010: oled_data = 16'b1011001001001001;
				18'b011010001000100010: oled_data = 16'b1011001001001001;
				18'b011010001010100010: oled_data = 16'b1011001001001001;
				18'b011010001100100010: oled_data = 16'b1010101000101000;
				18'b011010001110100010: oled_data = 16'b1011001001001001;
				18'b011010010000100010: oled_data = 16'b1001000101100110;
				18'b011010010010100010: oled_data = 16'b1000100101000110;
				18'b011010010100100010: oled_data = 16'b1010101000001001;
				18'b011010010110100010: oled_data = 16'b1011001001001001;
				18'b011010011000100010: oled_data = 16'b1011001001001001;
				18'b011010011010100010: oled_data = 16'b1011001001001001;
				18'b011010011100100010: oled_data = 16'b1011001001001001;
				18'b011010011110100010: oled_data = 16'b1011001001001001;
				18'b011010100000100010: oled_data = 16'b1011001000101001;
				18'b011010100010100010: oled_data = 16'b1011001000101000;
				18'b011010100100100010: oled_data = 16'b1010101000101000;
				18'b011010100110100010: oled_data = 16'b1010101000101000;
				18'b011000011000100011: oled_data = 16'b0110101010101100;
				18'b011000011010100011: oled_data = 16'b1010001110101111;
				18'b011000011100100011: oled_data = 16'b1101110011110100;
				18'b011000011110100011: oled_data = 16'b1101010010010100;
				18'b011000100000100011: oled_data = 16'b1100001111110010;
				18'b011000100010100011: oled_data = 16'b1110010011110110;
				18'b011000100100100011: oled_data = 16'b1100110000110011;
				18'b011000100110100011: oled_data = 16'b1011001101010000;
				18'b011000101000100011: oled_data = 16'b1100110000110100;
				18'b011000101010100011: oled_data = 16'b1101010100110101;
				18'b011000101100100011: oled_data = 16'b1010010011010010;
				18'b011000101110100011: oled_data = 16'b0011100110000101;
				18'b011000110000100011: oled_data = 16'b0101001001001000;
				18'b011000110010100011: oled_data = 16'b1101011001011000;
				18'b011000110100100011: oled_data = 16'b1110111011011010;
				18'b011000110110100011: oled_data = 16'b1101010101010101;
				18'b011000111000100011: oled_data = 16'b1101010010010100;
				18'b011000111010100011: oled_data = 16'b1101010010010101;
				18'b011000111100100011: oled_data = 16'b1101110011010110;
				18'b011000111110100011: oled_data = 16'b1101110011010101;
				18'b011001000000100011: oled_data = 16'b1110010011010101;
				18'b011001000010100011: oled_data = 16'b1101110011010101;
				18'b011001000100100011: oled_data = 16'b1101110011010110;
				18'b011001000110100011: oled_data = 16'b1101010011010101;
				18'b011001001000100011: oled_data = 16'b1110011001111001;
				18'b011001001010100011: oled_data = 16'b1110111100111100;
				18'b011001001100100011: oled_data = 16'b1101111000011001;
				18'b011001001110100011: oled_data = 16'b1100010010110100;
				18'b011001010000100011: oled_data = 16'b0111101100101100;
				18'b011001010010100011: oled_data = 16'b0011100101100101;
				18'b011001010100100011: oled_data = 16'b0100000110100110;
				18'b011001010110100011: oled_data = 16'b1001010000110000;
				18'b011001011000100011: oled_data = 16'b1101011000011000;
				18'b011001011010100011: oled_data = 16'b1100110100010101;
				18'b011001011100100011: oled_data = 16'b1100110011010101;
				18'b011001011110100011: oled_data = 16'b1110011010111010;
				18'b011001100000100011: oled_data = 16'b1110111100111011;
				18'b011001100010100011: oled_data = 16'b1110011001111010;
				18'b011001100100100011: oled_data = 16'b1011001110110001;
				18'b011001100110100011: oled_data = 16'b1011101111010010;
				18'b011001101000100011: oled_data = 16'b1100110001110100;
				18'b011001101010100011: oled_data = 16'b1101010001110100;
				18'b011001101100100011: oled_data = 16'b1101010001110101;
				18'b011001101110100011: oled_data = 16'b1101110010110101;
				18'b011001110000100011: oled_data = 16'b1101110011010110;
				18'b011001110010100011: oled_data = 16'b1101110011010110;
				18'b011001110100100011: oled_data = 16'b1101110011010110;
				18'b011001110110100011: oled_data = 16'b1101110010110101;
				18'b011001111000100011: oled_data = 16'b1101010010010101;
				18'b011001111010100011: oled_data = 16'b1101010001110100;
				18'b011001111100100011: oled_data = 16'b1101010001110011;
				18'b011001111110100011: oled_data = 16'b1110110100010100;
				18'b011010000000100011: oled_data = 16'b1011101100101100;
				18'b011010000010100011: oled_data = 16'b1011001000101001;
				18'b011010000100100011: oled_data = 16'b1011001001001001;
				18'b011010000110100011: oled_data = 16'b1011001001001001;
				18'b011010001000100011: oled_data = 16'b1011101001001001;
				18'b011010001010100011: oled_data = 16'b1011001000101001;
				18'b011010001100100011: oled_data = 16'b1010101000101001;
				18'b011010001110100011: oled_data = 16'b1010000111101000;
				18'b011010010000100011: oled_data = 16'b1000100101000110;
				18'b011010010010100011: oled_data = 16'b1001100111000111;
				18'b011010010100100011: oled_data = 16'b1011001001001001;
				18'b011010010110100011: oled_data = 16'b1011001001001001;
				18'b011010011000100011: oled_data = 16'b1011001001001001;
				18'b011010011010100011: oled_data = 16'b1011001001001001;
				18'b011010011100100011: oled_data = 16'b1011001000101001;
				18'b011010011110100011: oled_data = 16'b1011001001001001;
				18'b011010100000100011: oled_data = 16'b1011001000101001;
				18'b011010100010100011: oled_data = 16'b1011001000101000;
				18'b011010100100100011: oled_data = 16'b1010101000101000;
				18'b011010100110100011: oled_data = 16'b1010101000101000;
				18'b011000011000100100: oled_data = 16'b0011100111100111;
				18'b011000011010100100: oled_data = 16'b1010001110110000;
				18'b011000011100100100: oled_data = 16'b1110010011110110;
				18'b011000011110100100: oled_data = 16'b1101110011010101;
				18'b011000100000100100: oled_data = 16'b1011101111010001;
				18'b011000100010100100: oled_data = 16'b1100110001010011;
				18'b011000100100100100: oled_data = 16'b1100110001010100;
				18'b011000100110100100: oled_data = 16'b1011001101010000;
				18'b011000101000100100: oled_data = 16'b1011001110110001;
				18'b011000101010100100: oled_data = 16'b1101110011010101;
				18'b011000101100100100: oled_data = 16'b1110111010011010;
				18'b011000101110100100: oled_data = 16'b1011110110110101;
				18'b011000110000100100: oled_data = 16'b0100101000000111;
				18'b011000110010100100: oled_data = 16'b0110001011001010;
				18'b011000110100100100: oled_data = 16'b1101111010111010;
				18'b011000110110100100: oled_data = 16'b1110011010111001;
				18'b011000111000100100: oled_data = 16'b1100110100010101;
				18'b011000111010100100: oled_data = 16'b1101010001110100;
				18'b011000111100100100: oled_data = 16'b1101110011010101;
				18'b011000111110100100: oled_data = 16'b1101110011010101;
				18'b011001000000100100: oled_data = 16'b1101110011010101;
				18'b011001000010100100: oled_data = 16'b1101110011010101;
				18'b011001000100100100: oled_data = 16'b1101110011010101;
				18'b011001000110100100: oled_data = 16'b1101010011010101;
				18'b011001001000100100: oled_data = 16'b1110011001111001;
				18'b011001001010100100: oled_data = 16'b1110111100011011;
				18'b011001001100100100: oled_data = 16'b1001110001110001;
				18'b011001001110100100: oled_data = 16'b0100100111000111;
				18'b011001010000100100: oled_data = 16'b0011000100100100;
				18'b011001010010100100: oled_data = 16'b0110101011101100;
				18'b011001010100100100: oled_data = 16'b1100111000010111;
				18'b011001010110100100: oled_data = 16'b1111011101011100;
				18'b011001011000100100: oled_data = 16'b1110111100111011;
				18'b011001011010100100: oled_data = 16'b1110011010011010;
				18'b011001011100100100: oled_data = 16'b1101010101010110;
				18'b011001011110100100: oled_data = 16'b1101010110110111;
				18'b011001100000100100: oled_data = 16'b1110111100011011;
				18'b011001100010100100: oled_data = 16'b1110111100111011;
				18'b011001100100100100: oled_data = 16'b1100110101010110;
				18'b011001100110100100: oled_data = 16'b1011001110010000;
				18'b011001101000100100: oled_data = 16'b1101010010010100;
				18'b011001101010100100: oled_data = 16'b1101110011010110;
				18'b011001101100100100: oled_data = 16'b1101110011010110;
				18'b011001101110100100: oled_data = 16'b1101110011010110;
				18'b011001110000100100: oled_data = 16'b1101110011010101;
				18'b011001110010100100: oled_data = 16'b1101110011010101;
				18'b011001110100100100: oled_data = 16'b1101110011010101;
				18'b011001110110100100: oled_data = 16'b1101010001110100;
				18'b011001111000100100: oled_data = 16'b1101110010110101;
				18'b011001111010100100: oled_data = 16'b1101110011010101;
				18'b011001111100100100: oled_data = 16'b1101110010110011;
				18'b011001111110100100: oled_data = 16'b1110110011110100;
				18'b011010000000100100: oled_data = 16'b1011001010101011;
				18'b011010000010100100: oled_data = 16'b1011001000101001;
				18'b011010000100100100: oled_data = 16'b1011001001001001;
				18'b011010000110100100: oled_data = 16'b1011001001001001;
				18'b011010001000100100: oled_data = 16'b1011001001001001;
				18'b011010001010100100: oled_data = 16'b1010101000101000;
				18'b011010001100100100: oled_data = 16'b1011001000101001;
				18'b011010001110100100: oled_data = 16'b1001000101100110;
				18'b011010010000100100: oled_data = 16'b1001000101100111;
				18'b011010010010100100: oled_data = 16'b1011001000101001;
				18'b011010010100100100: oled_data = 16'b1011001001001001;
				18'b011010010110100100: oled_data = 16'b1011001000101001;
				18'b011010011000100100: oled_data = 16'b1011001001001001;
				18'b011010011010100100: oled_data = 16'b1011001001001001;
				18'b011010011100100100: oled_data = 16'b1011001001001001;
				18'b011010011110100100: oled_data = 16'b1011001001001001;
				18'b011010100000100100: oled_data = 16'b1011001000101001;
				18'b011010100010100100: oled_data = 16'b1011001000101000;
				18'b011010100100100100: oled_data = 16'b1010101000101000;
				18'b011010100110100100: oled_data = 16'b1010101000101000;
				18'b011000011000100101: oled_data = 16'b0011000111100111;
				18'b011000011010100101: oled_data = 16'b1001101101001111;
				18'b011000011100100101: oled_data = 16'b1101110011010101;
				18'b011000011110100101: oled_data = 16'b1101110011110110;
				18'b011000100000100101: oled_data = 16'b1100110001010011;
				18'b011000100010100101: oled_data = 16'b1011001110010001;
				18'b011000100100100101: oled_data = 16'b1101010001110100;
				18'b011000100110100101: oled_data = 16'b1011101110110001;
				18'b011000101000100101: oled_data = 16'b1011001111110010;
				18'b011000101010100101: oled_data = 16'b1101110011010101;
				18'b011000101100100101: oled_data = 16'b1110011000011000;
				18'b011000101110100101: oled_data = 16'b1111011101111011;
				18'b011000110000100101: oled_data = 16'b1100110111110110;
				18'b011000110010100101: oled_data = 16'b0100101000000111;
				18'b011000110100100101: oled_data = 16'b0111101101101101;
				18'b011000110110100101: oled_data = 16'b1110111100011010;
				18'b011000111000100101: oled_data = 16'b1101111001011000;
				18'b011000111010100101: oled_data = 16'b1100110011010100;
				18'b011000111100100101: oled_data = 16'b1101110010010100;
				18'b011000111110100101: oled_data = 16'b1101110011010101;
				18'b011001000000100101: oled_data = 16'b1110010011010101;
				18'b011001000010100101: oled_data = 16'b1101110011010101;
				18'b011001000100100101: oled_data = 16'b1101110011010101;
				18'b011001000110100101: oled_data = 16'b1101110011110110;
				18'b011001001000100101: oled_data = 16'b1100010110010110;
				18'b011001001010100101: oled_data = 16'b0110101100001100;
				18'b011001001100100101: oled_data = 16'b0011000100100101;
				18'b011001001110100101: oled_data = 16'b0100000111000111;
				18'b011001010000100101: oled_data = 16'b1001110001110001;
				18'b011001010010100101: oled_data = 16'b1110111100011011;
				18'b011001010100100101: oled_data = 16'b1110111100111100;
				18'b011001010110100101: oled_data = 16'b1110111100011011;
				18'b011001011000100101: oled_data = 16'b1110111100011010;
				18'b011001011010100101: oled_data = 16'b1110111100011011;
				18'b011001011100100101: oled_data = 16'b1110111100011011;
				18'b011001011110100101: oled_data = 16'b1101111010011001;
				18'b011001100000100101: oled_data = 16'b1110111100011010;
				18'b011001100010100101: oled_data = 16'b1110111100011010;
				18'b011001100100100101: oled_data = 16'b1110011011111010;
				18'b011001100110100101: oled_data = 16'b1011110001010010;
				18'b011001101000100101: oled_data = 16'b1100001111110010;
				18'b011001101010100101: oled_data = 16'b1101110010110101;
				18'b011001101100100101: oled_data = 16'b1101110011010110;
				18'b011001101110100101: oled_data = 16'b1101110011010101;
				18'b011001110000100101: oled_data = 16'b1101110011010101;
				18'b011001110010100101: oled_data = 16'b1101110011010110;
				18'b011001110100100101: oled_data = 16'b1101010010010100;
				18'b011001110110100101: oled_data = 16'b1101010010010100;
				18'b011001111000100101: oled_data = 16'b1101110011010110;
				18'b011001111010100101: oled_data = 16'b1101110010110101;
				18'b011001111100100101: oled_data = 16'b1101110010110100;
				18'b011001111110100101: oled_data = 16'b1110010011010011;
				18'b011010000000100101: oled_data = 16'b1010101001101001;
				18'b011010000010100101: oled_data = 16'b1011001001001001;
				18'b011010000100100101: oled_data = 16'b1011001001001001;
				18'b011010000110100101: oled_data = 16'b1011001001001001;
				18'b011010001000100101: oled_data = 16'b1011101010101010;
				18'b011010001010100101: oled_data = 16'b1011001010001001;
				18'b011010001100100101: oled_data = 16'b1010000111100111;
				18'b011010001110100101: oled_data = 16'b1000100101000110;
				18'b011010010000100101: oled_data = 16'b1010000111101001;
				18'b011010010010100101: oled_data = 16'b1011001001001001;
				18'b011010010100100101: oled_data = 16'b1011001000101001;
				18'b011010010110100101: oled_data = 16'b1011101110101111;
				18'b011010011000100101: oled_data = 16'b1011001010101011;
				18'b011010011010100101: oled_data = 16'b1011001001001001;
				18'b011010011100100101: oled_data = 16'b1011101010001010;
				18'b011010011110100101: oled_data = 16'b1011001001001001;
				18'b011010100000100101: oled_data = 16'b1011001000101001;
				18'b011010100010100101: oled_data = 16'b1011001000101000;
				18'b011010100100100101: oled_data = 16'b1010101000101000;
				18'b011010100110100101: oled_data = 16'b1010101000101000;
				18'b011000011000100110: oled_data = 16'b0100000111100111;
				18'b011000011010100110: oled_data = 16'b1011110000110010;
				18'b011000011100100110: oled_data = 16'b1101010001010100;
				18'b011000011110100110: oled_data = 16'b1101110011010110;
				18'b011000100000100110: oled_data = 16'b1101110010110101;
				18'b011000100010100110: oled_data = 16'b1100001111110010;
				18'b011000100100100110: oled_data = 16'b1011101110110001;
				18'b011000100110100110: oled_data = 16'b1011001101110001;
				18'b011000101000100110: oled_data = 16'b1011110000110011;
				18'b011000101010100110: oled_data = 16'b1110010111111000;
				18'b011000101100100110: oled_data = 16'b1101010110110111;
				18'b011000101110100110: oled_data = 16'b1110111100111011;
				18'b011000110000100110: oled_data = 16'b1111011101111100;
				18'b011000110010100110: oled_data = 16'b1100111000110111;
				18'b011000110100100110: oled_data = 16'b0100100111100111;
				18'b011000110110100110: oled_data = 16'b1001010001010000;
				18'b011000111000100110: oled_data = 16'b1110111101011011;
				18'b011000111010100110: oled_data = 16'b1101010111110111;
				18'b011000111100100110: oled_data = 16'b1101010010010100;
				18'b011000111110100110: oled_data = 16'b1101110010110101;
				18'b011001000000100110: oled_data = 16'b1110010011010101;
				18'b011001000010100110: oled_data = 16'b1101110011010101;
				18'b011001000100100110: oled_data = 16'b1110010011110110;
				18'b011001000110100110: oled_data = 16'b1100010000110011;
				18'b011001001000100110: oled_data = 16'b0101000111101000;
				18'b011001001010100110: oled_data = 16'b0011000110000101;
				18'b011001001100100110: oled_data = 16'b0111101110101110;
				18'b011001001110100110: oled_data = 16'b1011110101010101;
				18'b011001010000100110: oled_data = 16'b1101111000011000;
				18'b011001010010100110: oled_data = 16'b1110111100111011;
				18'b011001010100100110: oled_data = 16'b1110111100011010;
				18'b011001010110100110: oled_data = 16'b1110111100011010;
				18'b011001011000100110: oled_data = 16'b1110011100011010;
				18'b011001011010100110: oled_data = 16'b1110011100011010;
				18'b011001011100100110: oled_data = 16'b1110111100011010;
				18'b011001011110100110: oled_data = 16'b1110111100011011;
				18'b011001100000100110: oled_data = 16'b1110111100011010;
				18'b011001100010100110: oled_data = 16'b1110111100011010;
				18'b011001100100100110: oled_data = 16'b1110111100111010;
				18'b011001100110100110: oled_data = 16'b1101111001011000;
				18'b011001101000100110: oled_data = 16'b1011010000010001;
				18'b011001101010100110: oled_data = 16'b1101010001110100;
				18'b011001101100100110: oled_data = 16'b1101110011010101;
				18'b011001101110100110: oled_data = 16'b1101110011010101;
				18'b011001110000100110: oled_data = 16'b1101010010010100;
				18'b011001110010100110: oled_data = 16'b1101110010110101;
				18'b011001110100100110: oled_data = 16'b1101010010010101;
				18'b011001110110100110: oled_data = 16'b1101110011010101;
				18'b011001111000100110: oled_data = 16'b1101110011010101;
				18'b011001111010100110: oled_data = 16'b1101110010110101;
				18'b011001111100100110: oled_data = 16'b1101110011010100;
				18'b011001111110100110: oled_data = 16'b1101110001110001;
				18'b011010000000100110: oled_data = 16'b1010101000101000;
				18'b011010000010100110: oled_data = 16'b1011001001001001;
				18'b011010000100100110: oled_data = 16'b1011001010101010;
				18'b011010000110100110: oled_data = 16'b1101010000110001;
				18'b011010001000100110: oled_data = 16'b1110010010110011;
				18'b011010001010100110: oled_data = 16'b1100101110101111;
				18'b011010001100100110: oled_data = 16'b1010001000001000;
				18'b011010001110100110: oled_data = 16'b1001100110000111;
				18'b011010010000100110: oled_data = 16'b1011001001101010;
				18'b011010010010100110: oled_data = 16'b1011001001001001;
				18'b011010010100100110: oled_data = 16'b1011001001101010;
				18'b011010010110100110: oled_data = 16'b1100011000111001;
				18'b011010011000100110: oled_data = 16'b1011001111110000;
				18'b011010011010100110: oled_data = 16'b1011001000001001;
				18'b011010011100100110: oled_data = 16'b1011001000101001;
				18'b011010011110100110: oled_data = 16'b1011001000101001;
				18'b011010100000100110: oled_data = 16'b1011001000101001;
				18'b011010100010100110: oled_data = 16'b1011001000101000;
				18'b011010100100100110: oled_data = 16'b1010101000101000;
				18'b011010100110100110: oled_data = 16'b1010101000101000;
				18'b011000011000100111: oled_data = 16'b0100000110100111;
				18'b011000011010100111: oled_data = 16'b1101010010010100;
				18'b011000011100100111: oled_data = 16'b1101010010010100;
				18'b011000011110100111: oled_data = 16'b1101110011010101;
				18'b011000100000100111: oled_data = 16'b1110010011010110;
				18'b011000100010100111: oled_data = 16'b1100110000110011;
				18'b011000100100100111: oled_data = 16'b1011001101110000;
				18'b011000100110100111: oled_data = 16'b1010101100110000;
				18'b011000101000100111: oled_data = 16'b1100010001110100;
				18'b011000101010100111: oled_data = 16'b1111011100011011;
				18'b011000101100100111: oled_data = 16'b1101010111110111;
				18'b011000101110100111: oled_data = 16'b1101011001111000;
				18'b011000110000100111: oled_data = 16'b1100010111110110;
				18'b011000110010100111: oled_data = 16'b1010110100110100;
				18'b011000110100100111: oled_data = 16'b0110001011001010;
				18'b011000110110100111: oled_data = 16'b0100000110000110;
				18'b011000111000100111: oled_data = 16'b1101111001111000;
				18'b011000111010100111: oled_data = 16'b1110111100011010;
				18'b011000111100100111: oled_data = 16'b1101010111010111;
				18'b011000111110100111: oled_data = 16'b1100110010010100;
				18'b011001000000100111: oled_data = 16'b1101110010110101;
				18'b011001000010100111: oled_data = 16'b1101110011010101;
				18'b011001000100100111: oled_data = 16'b1110010011110110;
				18'b011001000110100111: oled_data = 16'b1000101011001101;
				18'b011001001000100111: oled_data = 16'b0011100100100101;
				18'b011001001010100111: oled_data = 16'b0101001010001001;
				18'b011001001100100111: oled_data = 16'b1100111000110111;
				18'b011001001110100111: oled_data = 16'b1101111001111001;
				18'b011001010000100111: oled_data = 16'b1101111000011000;
				18'b011001010010100111: oled_data = 16'b1110111101011011;
				18'b011001010100100111: oled_data = 16'b1110111100111011;
				18'b011001010110100111: oled_data = 16'b1110111100011011;
				18'b011001011000100111: oled_data = 16'b1110111100011010;
				18'b011001011010100111: oled_data = 16'b1110111100011010;
				18'b011001011100100111: oled_data = 16'b1110111100011010;
				18'b011001011110100111: oled_data = 16'b1110111100011010;
				18'b011001100000100111: oled_data = 16'b1110111100011010;
				18'b011001100010100111: oled_data = 16'b1110111100011010;
				18'b011001100100100111: oled_data = 16'b1110111100011010;
				18'b011001100110100111: oled_data = 16'b1110111100111011;
				18'b011001101000100111: oled_data = 16'b1101011000111000;
				18'b011001101010100111: oled_data = 16'b1011010000010010;
				18'b011001101100100111: oled_data = 16'b1101110010110101;
				18'b011001101110100111: oled_data = 16'b1101110011010110;
				18'b011001110000100111: oled_data = 16'b1101110010110101;
				18'b011001110010100111: oled_data = 16'b1100010000110011;
				18'b011001110100100111: oled_data = 16'b1101110011010101;
				18'b011001110110100111: oled_data = 16'b1101110011010101;
				18'b011001111000100111: oled_data = 16'b1101110011010101;
				18'b011001111010100111: oled_data = 16'b1101010010110101;
				18'b011001111100100111: oled_data = 16'b1101110011110100;
				18'b011001111110100111: oled_data = 16'b1101010000110000;
				18'b011010000000100111: oled_data = 16'b1010101000101000;
				18'b011010000010100111: oled_data = 16'b1011001001001001;
				18'b011010000100100111: oled_data = 16'b1101010001010001;
				18'b011010000110100111: oled_data = 16'b1110110011110011;
				18'b011010001000100111: oled_data = 16'b1100001100001100;
				18'b011010001010100111: oled_data = 16'b1011001000101001;
				18'b011010001100100111: oled_data = 16'b1011001001001001;
				18'b011010001110100111: oled_data = 16'b1011001001001001;
				18'b011010010000100111: oled_data = 16'b1011001001101010;
				18'b011010010010100111: oled_data = 16'b1011001000101001;
				18'b011010010100100111: oled_data = 16'b1011101111110000;
				18'b011010010110100111: oled_data = 16'b1100011100011100;
				18'b011010011000100111: oled_data = 16'b1011110111010111;
				18'b011010011010100111: oled_data = 16'b1011001001001001;
				18'b011010011100100111: oled_data = 16'b1011001001001001;
				18'b011010011110100111: oled_data = 16'b1011001000101001;
				18'b011010100000100111: oled_data = 16'b1010101000101000;
				18'b011010100010100111: oled_data = 16'b1010101000101000;
				18'b011010100100100111: oled_data = 16'b1010000111101000;
				18'b011010100110100111: oled_data = 16'b1010101000001000;
				18'b011000011000101000: oled_data = 16'b0110001000101000;
				18'b011000011010101000: oled_data = 16'b1101110010110101;
				18'b011000011100101000: oled_data = 16'b1101110011010110;
				18'b011000011110101000: oled_data = 16'b1101110011010110;
				18'b011000100000101000: oled_data = 16'b1101110011010110;
				18'b011000100010101000: oled_data = 16'b1101110010110101;
				18'b011000100100101000: oled_data = 16'b1011001101110000;
				18'b011000100110101000: oled_data = 16'b1011001101110000;
				18'b011000101000101000: oled_data = 16'b1100110011010101;
				18'b011000101010101000: oled_data = 16'b1010110100010011;
				18'b011000101100101000: oled_data = 16'b0101001001001000;
				18'b011000101110101000: oled_data = 16'b0011100110100110;
				18'b011000110000101000: oled_data = 16'b0011000101100101;
				18'b011000110010101000: oled_data = 16'b0011000101000100;
				18'b011000110100101000: oled_data = 16'b0100000110100110;
				18'b011000110110101000: oled_data = 16'b0110101011101011;
				18'b011000111000101000: oled_data = 16'b1101011001111000;
				18'b011000111010101000: oled_data = 16'b1110111100011010;
				18'b011000111100101000: oled_data = 16'b1110011011111010;
				18'b011000111110101000: oled_data = 16'b1101010110010111;
				18'b011001000000101000: oled_data = 16'b1100010001010011;
				18'b011001000010101000: oled_data = 16'b1101110010110101;
				18'b011001000100101000: oled_data = 16'b1110010011010110;
				18'b011001000110101000: oled_data = 16'b1011110000110010;
				18'b011001001000101000: oled_data = 16'b0110101010101010;
				18'b011001001010101000: oled_data = 16'b0011100110000110;
				18'b011001001100101000: oled_data = 16'b0011100101100101;
				18'b011001001110101000: oled_data = 16'b0101001001001000;
				18'b011001010000101000: oled_data = 16'b0111101101101101;
				18'b011001010010101000: oled_data = 16'b1010010011110011;
				18'b011001010100101000: oled_data = 16'b1100111000010111;
				18'b011001010110101000: oled_data = 16'b1101111010111010;
				18'b011001011000101000: oled_data = 16'b1110111100111011;
				18'b011001011010101000: oled_data = 16'b1110111101011011;
				18'b011001011100101000: oled_data = 16'b1110111100011011;
				18'b011001011110101000: oled_data = 16'b1110111100011010;
				18'b011001100000101000: oled_data = 16'b1110111100011010;
				18'b011001100010101000: oled_data = 16'b1110111100011010;
				18'b011001100100101000: oled_data = 16'b1110111100011010;
				18'b011001100110101000: oled_data = 16'b1110011100011010;
				18'b011001101000101000: oled_data = 16'b1110111100111010;
				18'b011001101010101000: oled_data = 16'b1100110110110110;
				18'b011001101100101000: oled_data = 16'b1100010001110011;
				18'b011001101110101000: oled_data = 16'b1101110011110110;
				18'b011001110000101000: oled_data = 16'b1101010001110100;
				18'b011001110010101000: oled_data = 16'b1101010010010100;
				18'b011001110100101000: oled_data = 16'b1101010001110100;
				18'b011001110110101000: oled_data = 16'b1101110011010101;
				18'b011001111000101000: oled_data = 16'b1101110011010101;
				18'b011001111010101000: oled_data = 16'b1101110010110101;
				18'b011001111100101000: oled_data = 16'b1101110011110100;
				18'b011001111110101000: oled_data = 16'b1100101111001111;
				18'b011010000000101000: oled_data = 16'b1010101000001000;
				18'b011010000010101000: oled_data = 16'b1011101011101100;
				18'b011010000100101000: oled_data = 16'b1110010011110100;
				18'b011010000110101000: oled_data = 16'b1100101101101110;
				18'b011010001000101000: oled_data = 16'b1011001000101001;
				18'b011010001010101000: oled_data = 16'b1011001001001001;
				18'b011010001100101000: oled_data = 16'b1011001001001001;
				18'b011010001110101000: oled_data = 16'b1011001001001001;
				18'b011010010000101000: oled_data = 16'b1011001001001001;
				18'b011010010010101000: oled_data = 16'b1011001001001001;
				18'b011010010100101000: oled_data = 16'b1100010110010110;
				18'b011010010110101000: oled_data = 16'b1011111100011100;
				18'b011010011000101000: oled_data = 16'b1011111011111011;
				18'b011010011010101000: oled_data = 16'b1011001101101110;
				18'b011010011100101000: oled_data = 16'b1011001000001000;
				18'b011010011110101000: oled_data = 16'b1010101000001000;
				18'b011010100000101000: oled_data = 16'b1010001000001000;
				18'b011010100010101000: oled_data = 16'b1010001000001000;
				18'b011010100100101000: oled_data = 16'b1010101000001000;
				18'b011010100110101000: oled_data = 16'b1010101000001000;
				18'b011000011000101001: oled_data = 16'b1000101110001101;
				18'b011000011010101001: oled_data = 16'b1101110010110110;
				18'b011000011100101001: oled_data = 16'b1101110011010110;
				18'b011000011110101001: oled_data = 16'b1101110011010110;
				18'b011000100000101001: oled_data = 16'b1101110011010110;
				18'b011000100010101001: oled_data = 16'b1101110011010110;
				18'b011000100100101001: oled_data = 16'b1011101110110001;
				18'b011000100110101001: oled_data = 16'b1011001101110001;
				18'b011000101000101001: oled_data = 16'b1100110100010110;
				18'b011000101010101001: oled_data = 16'b1001110010010001;
				18'b011000101100101001: oled_data = 16'b0110101100001100;
				18'b011000101110101001: oled_data = 16'b1000001111001111;
				18'b011000110000101001: oled_data = 16'b1010010010110010;
				18'b011000110010101001: oled_data = 16'b1011010110010101;
				18'b011000110100101001: oled_data = 16'b1101011001011000;
				18'b011000110110101001: oled_data = 16'b1110111100111011;
				18'b011000111000101001: oled_data = 16'b1110011100011010;
				18'b011000111010101001: oled_data = 16'b1110011011111010;
				18'b011000111100101001: oled_data = 16'b1110011100011010;
				18'b011000111110101001: oled_data = 16'b1110111100011011;
				18'b011001000000101001: oled_data = 16'b1101010111010111;
				18'b011001000010101001: oled_data = 16'b1100010010010011;
				18'b011001000100101001: oled_data = 16'b1101110011010101;
				18'b011001000110101001: oled_data = 16'b1101010100010101;
				18'b011001001000101001: oled_data = 16'b1110011010011010;
				18'b011001001010101001: oled_data = 16'b1100010110110110;
				18'b011001001100101001: oled_data = 16'b1000101111101111;
				18'b011001001110101001: oled_data = 16'b0101101010001010;
				18'b011001010000101001: oled_data = 16'b0100000110100110;
				18'b011001010010101001: oled_data = 16'b0011100101000101;
				18'b011001010100101001: oled_data = 16'b0011100110000101;
				18'b011001010110101001: oled_data = 16'b0100101000101000;
				18'b011001011000101001: oled_data = 16'b0110101100001011;
				18'b011001011010101001: oled_data = 16'b1000110000101111;
				18'b011001011100101001: oled_data = 16'b1101011001011000;
				18'b011001011110101001: oled_data = 16'b1110111100011011;
				18'b011001100000101001: oled_data = 16'b1110111100011010;
				18'b011001100010101001: oled_data = 16'b1110111100011010;
				18'b011001100100101001: oled_data = 16'b1110111100011010;
				18'b011001100110101001: oled_data = 16'b1110011100011010;
				18'b011001101000101001: oled_data = 16'b1110011100011010;
				18'b011001101010101001: oled_data = 16'b1111011101011100;
				18'b011001101100101001: oled_data = 16'b1011110011110011;
				18'b011001101110101001: oled_data = 16'b1100010000110011;
				18'b011001110000101001: oled_data = 16'b1101010010010100;
				18'b011001110010101001: oled_data = 16'b1101110011010101;
				18'b011001110100101001: oled_data = 16'b1101010010110101;
				18'b011001110110101001: oled_data = 16'b1101010001110100;
				18'b011001111000101001: oled_data = 16'b1101110010110101;
				18'b011001111010101001: oled_data = 16'b1101110010110101;
				18'b011001111100101001: oled_data = 16'b1101110011110100;
				18'b011001111110101001: oled_data = 16'b1100101110001110;
				18'b011010000000101001: oled_data = 16'b1011001000001000;
				18'b011010000010101001: oled_data = 16'b1100101110101110;
				18'b011010000100101001: oled_data = 16'b1110010010110010;
				18'b011010000110101001: oled_data = 16'b1011101010001010;
				18'b011010001000101001: oled_data = 16'b1011001001001001;
				18'b011010001010101001: oled_data = 16'b1011001001001001;
				18'b011010001100101001: oled_data = 16'b1011001001001001;
				18'b011010001110101001: oled_data = 16'b1011001001001001;
				18'b011010010000101001: oled_data = 16'b1011001000101001;
				18'b011010010010101001: oled_data = 16'b1011001101101110;
				18'b011010010100101001: oled_data = 16'b1100011011011011;
				18'b011010010110101001: oled_data = 16'b1011111011111011;
				18'b011010011000101001: oled_data = 16'b1011111100011100;
				18'b011010011010101001: oled_data = 16'b1011110101010101;
				18'b011010011100101001: oled_data = 16'b1010101000101000;
				18'b011010011110101001: oled_data = 16'b1011001000101000;
				18'b011010100000101001: oled_data = 16'b1011001000101000;
				18'b011010100010101001: oled_data = 16'b1010101000101000;
				18'b011010100100101001: oled_data = 16'b1010101000001000;
				18'b011010100110101001: oled_data = 16'b1010101000001000;
				18'b011000011000101010: oled_data = 16'b1010101111110000;
				18'b011000011010101010: oled_data = 16'b1110010010110110;
				18'b011000011100101010: oled_data = 16'b1101110011010110;
				18'b011000011110101010: oled_data = 16'b1101110011010110;
				18'b011000100000101010: oled_data = 16'b1101110011010110;
				18'b011000100010101010: oled_data = 16'b1101110010110101;
				18'b011000100100101010: oled_data = 16'b1011001110010001;
				18'b011000100110101010: oled_data = 16'b1011001101110001;
				18'b011000101000101010: oled_data = 16'b1101010110010111;
				18'b011000101010101010: oled_data = 16'b1110111100111011;
				18'b011000101100101010: oled_data = 16'b1110111100111011;
				18'b011000101110101010: oled_data = 16'b1111011100111011;
				18'b011000110000101010: oled_data = 16'b1110111100111011;
				18'b011000110010101010: oled_data = 16'b1110111100111011;
				18'b011000110100101010: oled_data = 16'b1110111100011011;
				18'b011000110110101010: oled_data = 16'b1110111011111010;
				18'b011000111000101010: oled_data = 16'b1110111011111010;
				18'b011000111010101010: oled_data = 16'b1110111011111010;
				18'b011000111100101010: oled_data = 16'b1110111100011010;
				18'b011000111110101010: oled_data = 16'b1110111100011010;
				18'b011001000000101010: oled_data = 16'b1110111100011010;
				18'b011001000010101010: oled_data = 16'b1101111001011000;
				18'b011001000100101010: oled_data = 16'b1100010100110100;
				18'b011001000110101010: oled_data = 16'b1101010101010101;
				18'b011001001000101010: oled_data = 16'b1110011011111010;
				18'b011001001010101010: oled_data = 16'b1110111100111011;
				18'b011001001100101010: oled_data = 16'b1110111100111011;
				18'b011001001110101010: oled_data = 16'b1110011011111010;
				18'b011001010000101010: oled_data = 16'b1101011000111000;
				18'b011001010010101010: oled_data = 16'b1011010100110100;
				18'b011001010100101010: oled_data = 16'b1001010001110001;
				18'b011001010110101010: oled_data = 16'b0111001100101100;
				18'b011001011000101010: oled_data = 16'b0110001011001011;
				18'b011001011010101010: oled_data = 16'b0101001001001000;
				18'b011001011100101010: oled_data = 16'b1011110110110101;
				18'b011001011110101010: oled_data = 16'b1110111100111011;
				18'b011001100000101010: oled_data = 16'b1110111100011010;
				18'b011001100010101010: oled_data = 16'b1110111100011010;
				18'b011001100100101010: oled_data = 16'b1110111100011010;
				18'b011001100110101010: oled_data = 16'b1110011100011010;
				18'b011001101000101010: oled_data = 16'b1110111100011010;
				18'b011001101010101010: oled_data = 16'b1101111000110111;
				18'b011001101100101010: oled_data = 16'b1101010100110100;
				18'b011001101110101010: oled_data = 16'b1100110010110011;
				18'b011001110000101010: oled_data = 16'b1101010010110100;
				18'b011001110010101010: oled_data = 16'b1101110010110101;
				18'b011001110100101010: oled_data = 16'b1101110010110101;
				18'b011001110110101010: oled_data = 16'b1101110010110101;
				18'b011001111000101010: oled_data = 16'b1101010010010100;
				18'b011001111010101010: oled_data = 16'b1100110001010100;
				18'b011001111100101010: oled_data = 16'b1101110011010100;
				18'b011001111110101010: oled_data = 16'b1100001101001101;
				18'b011010000000101010: oled_data = 16'b1010101000001000;
				18'b011010000010101010: oled_data = 16'b1101010000110000;
				18'b011010000100101010: oled_data = 16'b1101110000010000;
				18'b011010000110101010: oled_data = 16'b1011001001001001;
				18'b011010001000101010: oled_data = 16'b1011101001001001;
				18'b011010001010101010: oled_data = 16'b1011001001001001;
				18'b011010001100101010: oled_data = 16'b1011001001001001;
				18'b011010001110101010: oled_data = 16'b1011001001001001;
				18'b011010010000101010: oled_data = 16'b1011001000101001;
				18'b011010010010101010: oled_data = 16'b1011110101110101;
				18'b011010010100101010: oled_data = 16'b1011111100011100;
				18'b011010010110101010: oled_data = 16'b1011111011111011;
				18'b011010011000101010: oled_data = 16'b1011111011111100;
				18'b011010011010101010: oled_data = 16'b1100011010111010;
				18'b011010011100101010: oled_data = 16'b1011001100001100;
				18'b011010011110101010: oled_data = 16'b1010101000101000;
				18'b011010100000101010: oled_data = 16'b1011001000101001;
				18'b011010100010101010: oled_data = 16'b1010101000101000;
				18'b011010100100101010: oled_data = 16'b1010101000001000;
				18'b011010100110101010: oled_data = 16'b1010101000001000;
				18'b011000011000101011: oled_data = 16'b1011010000010001;
				18'b011000011010101011: oled_data = 16'b1110010010110110;
				18'b011000011100101011: oled_data = 16'b1101110011010110;
				18'b011000011110101011: oled_data = 16'b1101110011010110;
				18'b011000100000101011: oled_data = 16'b1101110011010110;
				18'b011000100010101011: oled_data = 16'b1101010010010101;
				18'b011000100100101011: oled_data = 16'b1011001101110000;
				18'b011000100110101011: oled_data = 16'b1011001101110001;
				18'b011000101000101011: oled_data = 16'b1101111000011000;
				18'b011000101010101011: oled_data = 16'b1110111100011010;
				18'b011000101100101011: oled_data = 16'b1110011100011010;
				18'b011000101110101011: oled_data = 16'b1110011100011010;
				18'b011000110000101011: oled_data = 16'b1110011100011010;
				18'b011000110010101011: oled_data = 16'b1110011011111010;
				18'b011000110100101011: oled_data = 16'b1110011100011010;
				18'b011000110110101011: oled_data = 16'b1110011011111010;
				18'b011000111000101011: oled_data = 16'b1110011011111010;
				18'b011000111010101011: oled_data = 16'b1110011011111010;
				18'b011000111100101011: oled_data = 16'b1110111100011010;
				18'b011000111110101011: oled_data = 16'b1110011100011010;
				18'b011001000000101011: oled_data = 16'b1110111011111010;
				18'b011001000010101011: oled_data = 16'b1110111100011010;
				18'b011001000100101011: oled_data = 16'b1110011010111001;
				18'b011001000110101011: oled_data = 16'b1101010111110111;
				18'b011001001000101011: oled_data = 16'b1110111100011010;
				18'b011001001010101011: oled_data = 16'b1110111100011010;
				18'b011001001100101011: oled_data = 16'b1110111100011010;
				18'b011001001110101011: oled_data = 16'b1110111100011010;
				18'b011001010000101011: oled_data = 16'b1110111100011011;
				18'b011001010010101011: oled_data = 16'b1110111100011011;
				18'b011001010100101011: oled_data = 16'b1111011100111100;
				18'b011001010110101011: oled_data = 16'b1110111100111100;
				18'b011001011000101011: oled_data = 16'b1110111011111011;
				18'b011001011010101011: oled_data = 16'b1110011011011010;
				18'b011001011100101011: oled_data = 16'b1110011011111010;
				18'b011001011110101011: oled_data = 16'b1110111100011010;
				18'b011001100000101011: oled_data = 16'b1110111100011010;
				18'b011001100010101011: oled_data = 16'b1110111100011010;
				18'b011001100100101011: oled_data = 16'b1110111100011010;
				18'b011001100110101011: oled_data = 16'b1110111100111011;
				18'b011001101000101011: oled_data = 16'b1101111001011000;
				18'b011001101010101011: oled_data = 16'b1101010100010100;
				18'b011001101100101011: oled_data = 16'b1110010101010101;
				18'b011001101110101011: oled_data = 16'b1101110101010101;
				18'b011001110000101011: oled_data = 16'b1101010011110100;
				18'b011001110010101011: oled_data = 16'b1100110011010100;
				18'b011001110100101011: oled_data = 16'b1101010010110100;
				18'b011001110110101011: oled_data = 16'b1101110011010101;
				18'b011001111000101011: oled_data = 16'b1110010011110110;
				18'b011001111010101011: oled_data = 16'b1101110010110101;
				18'b011001111100101011: oled_data = 16'b1101010010110011;
				18'b011001111110101011: oled_data = 16'b1011101100101101;
				18'b011010000000101011: oled_data = 16'b1011001000101001;
				18'b011010000010101011: oled_data = 16'b1101110001110001;
				18'b011010000100101011: oled_data = 16'b1100101101101110;
				18'b011010000110101011: oled_data = 16'b1011101000101001;
				18'b011010001000101011: oled_data = 16'b1011101001001001;
				18'b011010001010101011: oled_data = 16'b1011001001001001;
				18'b011010001100101011: oled_data = 16'b1011001001001001;
				18'b011010001110101011: oled_data = 16'b1011001000101001;
				18'b011010010000101011: oled_data = 16'b1010101011001011;
				18'b011010010010101011: oled_data = 16'b1011111010111010;
				18'b011010010100101011: oled_data = 16'b1011111011111011;
				18'b011010010110101011: oled_data = 16'b1011111011111011;
				18'b011010011000101011: oled_data = 16'b1011111011111100;
				18'b011010011010101011: oled_data = 16'b1100011100111100;
				18'b011010011100101011: oled_data = 16'b1011110011010011;
				18'b011010011110101011: oled_data = 16'b1010101000001000;
				18'b011010100000101011: oled_data = 16'b1011001000101001;
				18'b011010100010101011: oled_data = 16'b1010101000001000;
				18'b011010100100101011: oled_data = 16'b1010101000001000;
				18'b011010100110101011: oled_data = 16'b1010101000001000;
				18'b011000011000101100: oled_data = 16'b1011110001110010;
				18'b011000011010101100: oled_data = 16'b1101110011010110;
				18'b011000011100101100: oled_data = 16'b1101110010110101;
				18'b011000011110101100: oled_data = 16'b1101110010110101;
				18'b011000100000101100: oled_data = 16'b1101110011010110;
				18'b011000100010101100: oled_data = 16'b1100110001010100;
				18'b011000100100101100: oled_data = 16'b1011001101110000;
				18'b011000100110101100: oled_data = 16'b1011001110010001;
				18'b011000101000101100: oled_data = 16'b1101110111010111;
				18'b011000101010101100: oled_data = 16'b1110111100111010;
				18'b011000101100101100: oled_data = 16'b1110011100011010;
				18'b011000101110101100: oled_data = 16'b1110011011111010;
				18'b011000110000101100: oled_data = 16'b1110011011111010;
				18'b011000110010101100: oled_data = 16'b1110011011111010;
				18'b011000110100101100: oled_data = 16'b1110011011111010;
				18'b011000110110101100: oled_data = 16'b1110011011111010;
				18'b011000111000101100: oled_data = 16'b1110011011111010;
				18'b011000111010101100: oled_data = 16'b1110011100011010;
				18'b011000111100101100: oled_data = 16'b1110011100011010;
				18'b011000111110101100: oled_data = 16'b1110011100011010;
				18'b011001000000101100: oled_data = 16'b1110011100011010;
				18'b011001000010101100: oled_data = 16'b1110111100011010;
				18'b011001000100101100: oled_data = 16'b1110111100011010;
				18'b011001000110101100: oled_data = 16'b1110111100011010;
				18'b011001001000101100: oled_data = 16'b1110111100011010;
				18'b011001001010101100: oled_data = 16'b1110111100011010;
				18'b011001001100101100: oled_data = 16'b1110111100011010;
				18'b011001001110101100: oled_data = 16'b1110111100011010;
				18'b011001010000101100: oled_data = 16'b1110111100011010;
				18'b011001010010101100: oled_data = 16'b1110111100011010;
				18'b011001010100101100: oled_data = 16'b1110111100011010;
				18'b011001010110101100: oled_data = 16'b1110111100011011;
				18'b011001011000101100: oled_data = 16'b1110111100011010;
				18'b011001011010101100: oled_data = 16'b1110111100011011;
				18'b011001011100101100: oled_data = 16'b1110111100011010;
				18'b011001011110101100: oled_data = 16'b1110111100011010;
				18'b011001100000101100: oled_data = 16'b1110111100011010;
				18'b011001100010101100: oled_data = 16'b1110111100011010;
				18'b011001100100101100: oled_data = 16'b1110111100011010;
				18'b011001100110101100: oled_data = 16'b1101111000110111;
				18'b011001101000101100: oled_data = 16'b1101010101010101;
				18'b011001101010101100: oled_data = 16'b1101110100110101;
				18'b011001101100101100: oled_data = 16'b1101110101010101;
				18'b011001101110101100: oled_data = 16'b1101110101010101;
				18'b011001110000101100: oled_data = 16'b1101010110010110;
				18'b011001110010101100: oled_data = 16'b1110011011011010;
				18'b011001110100101100: oled_data = 16'b1101011000010111;
				18'b011001110110101100: oled_data = 16'b1100010100110100;
				18'b011001111000101100: oled_data = 16'b1101010011110101;
				18'b011001111010101100: oled_data = 16'b1101110011110101;
				18'b011001111100101100: oled_data = 16'b1101010010110100;
				18'b011001111110101100: oled_data = 16'b1011101100001100;
				18'b011010000000101100: oled_data = 16'b1011001001001001;
				18'b011010000010101100: oled_data = 16'b1101110010010010;
				18'b011010000100101100: oled_data = 16'b1100001011101100;
				18'b011010000110101100: oled_data = 16'b1011001000101001;
				18'b011010001000101100: oled_data = 16'b1011001001001001;
				18'b011010001010101100: oled_data = 16'b1011001001001001;
				18'b011010001100101100: oled_data = 16'b1011001001001001;
				18'b011010001110101100: oled_data = 16'b1011001000101001;
				18'b011010010000101100: oled_data = 16'b1011110000110001;
				18'b011010010010101100: oled_data = 16'b1011111100011100;
				18'b011010010100101100: oled_data = 16'b1011111011111011;
				18'b011010010110101100: oled_data = 16'b1011111011111011;
				18'b011010011000101100: oled_data = 16'b1011111011111011;
				18'b011010011010101100: oled_data = 16'b1100111100111101;
				18'b011010011100101100: oled_data = 16'b1011111000111000;
				18'b011010011110101100: oled_data = 16'b1010101010001010;
				18'b011010100000101100: oled_data = 16'b1010101000101000;
				18'b011010100010101100: oled_data = 16'b1010101000001000;
				18'b011010100100101100: oled_data = 16'b1010101000001000;
				18'b011010100110101100: oled_data = 16'b1010101000001000;
				18'b011000011000101101: oled_data = 16'b1011110001010010;
				18'b011000011010101101: oled_data = 16'b1101110011010101;
				18'b011000011100101101: oled_data = 16'b1101110010110101;
				18'b011000011110101101: oled_data = 16'b1101110010110101;
				18'b011000100000101101: oled_data = 16'b1101110011010110;
				18'b011000100010101101: oled_data = 16'b1100110000010011;
				18'b011000100100101101: oled_data = 16'b1011001101010000;
				18'b011000100110101101: oled_data = 16'b1011001101110000;
				18'b011000101000101101: oled_data = 16'b1011110000110010;
				18'b011000101010101101: oled_data = 16'b1110011011011010;
				18'b011000101100101101: oled_data = 16'b1110111100011010;
				18'b011000101110101101: oled_data = 16'b1110011011111010;
				18'b011000110000101101: oled_data = 16'b1110011011111010;
				18'b011000110010101101: oled_data = 16'b1110011011111010;
				18'b011000110100101101: oled_data = 16'b1110011011111010;
				18'b011000110110101101: oled_data = 16'b1110011011111010;
				18'b011000111000101101: oled_data = 16'b1110011011111010;
				18'b011000111010101101: oled_data = 16'b1110011011111010;
				18'b011000111100101101: oled_data = 16'b1110011011111010;
				18'b011000111110101101: oled_data = 16'b1110011011111010;
				18'b011001000000101101: oled_data = 16'b1110011011111010;
				18'b011001000010101101: oled_data = 16'b1110011011111010;
				18'b011001000100101101: oled_data = 16'b1110111011111010;
				18'b011001000110101101: oled_data = 16'b1110111100011010;
				18'b011001001000101101: oled_data = 16'b1110111011111010;
				18'b011001001010101101: oled_data = 16'b1110111011111010;
				18'b011001001100101101: oled_data = 16'b1110111011111010;
				18'b011001001110101101: oled_data = 16'b1110111100011010;
				18'b011001010000101101: oled_data = 16'b1110111100011010;
				18'b011001010010101101: oled_data = 16'b1110111100011010;
				18'b011001010100101101: oled_data = 16'b1110111100011010;
				18'b011001010110101101: oled_data = 16'b1110111100011010;
				18'b011001011000101101: oled_data = 16'b1110111100011010;
				18'b011001011010101101: oled_data = 16'b1110111100011010;
				18'b011001011100101101: oled_data = 16'b1110111100011010;
				18'b011001011110101101: oled_data = 16'b1110111100011010;
				18'b011001100000101101: oled_data = 16'b1110111100011010;
				18'b011001100010101101: oled_data = 16'b1110111100011010;
				18'b011001100100101101: oled_data = 16'b1101110111110111;
				18'b011001100110101101: oled_data = 16'b1101010100110101;
				18'b011001101000101101: oled_data = 16'b1101010100010101;
				18'b011001101010101101: oled_data = 16'b1101110101010101;
				18'b011001101100101101: oled_data = 16'b1101110101010110;
				18'b011001101110101101: oled_data = 16'b1101010100110101;
				18'b011001110000101101: oled_data = 16'b1101111001111000;
				18'b011001110010101101: oled_data = 16'b1110111100011010;
				18'b011001110100101101: oled_data = 16'b1101111011011001;
				18'b011001110110101101: oled_data = 16'b1110011010111001;
				18'b011001111000101101: oled_data = 16'b1110011001111001;
				18'b011001111010101101: oled_data = 16'b1101011000011000;
				18'b011001111100101101: oled_data = 16'b1100110100110101;
				18'b011001111110101101: oled_data = 16'b1011101011101100;
				18'b011010000000101101: oled_data = 16'b1011001001001010;
				18'b011010000010101101: oled_data = 16'b1101110001010001;
				18'b011010000100101101: oled_data = 16'b1011101010101011;
				18'b011010000110101101: oled_data = 16'b1011001000101001;
				18'b011010001000101101: oled_data = 16'b1011001001001001;
				18'b011010001010101101: oled_data = 16'b1011001001001001;
				18'b011010001100101101: oled_data = 16'b1011001001001001;
				18'b011010001110101101: oled_data = 16'b1011001001001001;
				18'b011010010000101101: oled_data = 16'b1100010110010111;
				18'b011010010010101101: oled_data = 16'b1011111100011100;
				18'b011010010100101101: oled_data = 16'b1011111011111011;
				18'b011010010110101101: oled_data = 16'b1011111011111011;
				18'b011010011000101101: oled_data = 16'b1011111011111011;
				18'b011010011010101101: oled_data = 16'b1100111100011100;
				18'b011010011100101101: oled_data = 16'b1011111011011011;
				18'b011010011110101101: oled_data = 16'b1010101101101101;
				18'b011010100000101101: oled_data = 16'b1010101000001000;
				18'b011010100010101101: oled_data = 16'b1010101000001000;
				18'b011010100100101101: oled_data = 16'b1010101000001000;
				18'b011010100110101101: oled_data = 16'b1010101000001000;
				18'b011000011000101110: oled_data = 16'b1011001111110001;
				18'b011000011010101110: oled_data = 16'b1101110011010101;
				18'b011000011100101110: oled_data = 16'b1101110010110101;
				18'b011000011110101110: oled_data = 16'b1101110010110101;
				18'b011000100000101110: oled_data = 16'b1101110011010101;
				18'b011000100010101110: oled_data = 16'b1100001111110010;
				18'b011000100100101110: oled_data = 16'b1011001101010000;
				18'b011000100110101110: oled_data = 16'b1011001101110000;
				18'b011000101000101110: oled_data = 16'b1011001101010000;
				18'b011000101010101110: oled_data = 16'b1011110001110011;
				18'b011000101100101110: oled_data = 16'b1110011010111010;
				18'b011000101110101110: oled_data = 16'b1110111100011010;
				18'b011000110000101110: oled_data = 16'b1110011011111010;
				18'b011000110010101110: oled_data = 16'b1110011011111010;
				18'b011000110100101110: oled_data = 16'b1110011011111010;
				18'b011000110110101110: oled_data = 16'b1110011011111010;
				18'b011000111000101110: oled_data = 16'b1110011011111010;
				18'b011000111010101110: oled_data = 16'b1110011011111010;
				18'b011000111100101110: oled_data = 16'b1110011011111010;
				18'b011000111110101110: oled_data = 16'b1110011011111010;
				18'b011001000000101110: oled_data = 16'b1110011011111010;
				18'b011001000010101110: oled_data = 16'b1110011011111010;
				18'b011001000100101110: oled_data = 16'b1110011011111010;
				18'b011001000110101110: oled_data = 16'b1110011011111010;
				18'b011001001000101110: oled_data = 16'b1110011011111010;
				18'b011001001010101110: oled_data = 16'b1110011011111010;
				18'b011001001100101110: oled_data = 16'b1110011011111010;
				18'b011001001110101110: oled_data = 16'b1110011011111010;
				18'b011001010000101110: oled_data = 16'b1110011011111010;
				18'b011001010010101110: oled_data = 16'b1110011011111010;
				18'b011001010100101110: oled_data = 16'b1110011011111010;
				18'b011001010110101110: oled_data = 16'b1110011011111010;
				18'b011001011000101110: oled_data = 16'b1110011100011010;
				18'b011001011010101110: oled_data = 16'b1110011100011010;
				18'b011001011100101110: oled_data = 16'b1110111100011010;
				18'b011001011110101110: oled_data = 16'b1110111100111010;
				18'b011001100000101110: oled_data = 16'b1110011011011001;
				18'b011001100010101110: oled_data = 16'b1100010100110100;
				18'b011001100100101110: oled_data = 16'b1101010100010100;
				18'b011001100110101110: oled_data = 16'b1101010100010100;
				18'b011001101000101110: oled_data = 16'b1101010011110100;
				18'b011001101010101110: oled_data = 16'b1101110100110101;
				18'b011001101100101110: oled_data = 16'b1101110100110101;
				18'b011001101110101110: oled_data = 16'b1101010110110110;
				18'b011001110000101110: oled_data = 16'b1110011100011010;
				18'b011001110010101110: oled_data = 16'b1110011011111010;
				18'b011001110100101110: oled_data = 16'b1101111010011001;
				18'b011001110110101110: oled_data = 16'b1110111100011010;
				18'b011001111000101110: oled_data = 16'b1110111100011010;
				18'b011001111010101110: oled_data = 16'b1110011100011010;
				18'b011001111100101110: oled_data = 16'b1101011000110111;
				18'b011001111110101110: oled_data = 16'b1011001011001011;
				18'b011010000000101110: oled_data = 16'b1011001001101010;
				18'b011010000010101110: oled_data = 16'b1101010000110000;
				18'b011010000100101110: oled_data = 16'b1011001001101010;
				18'b011010000110101110: oled_data = 16'b1011001000101001;
				18'b011010001000101110: oled_data = 16'b1011001000101001;
				18'b011010001010101110: oled_data = 16'b1011001000101001;
				18'b011010001100101110: oled_data = 16'b1011001000101001;
				18'b011010001110101110: oled_data = 16'b1011001010001010;
				18'b011010010000101110: oled_data = 16'b1100011001011001;
				18'b011010010010101110: oled_data = 16'b1011111011111100;
				18'b011010010100101110: oled_data = 16'b1011111011011011;
				18'b011010010110101110: oled_data = 16'b1011111011011011;
				18'b011010011000101110: oled_data = 16'b1011111011111011;
				18'b011010011010101110: oled_data = 16'b1100111100011100;
				18'b011010011100101110: oled_data = 16'b1011111100011100;
				18'b011010011110101110: oled_data = 16'b1011010010110010;
				18'b011010100000101110: oled_data = 16'b1010101000001000;
				18'b011010100010101110: oled_data = 16'b1010101000001000;
				18'b011010100100101110: oled_data = 16'b1010101000001000;
				18'b011010100110101110: oled_data = 16'b1010100111101000;
				18'b011000011000101111: oled_data = 16'b1011001111110001;
				18'b011000011010101111: oled_data = 16'b1101110010110101;
				18'b011000011100101111: oled_data = 16'b1101010001110100;
				18'b011000011110101111: oled_data = 16'b1101010001110100;
				18'b011000100000101111: oled_data = 16'b1101110010110101;
				18'b011000100010101111: oled_data = 16'b1011101111010010;
				18'b011000100100101111: oled_data = 16'b1011001101010000;
				18'b011000100110101111: oled_data = 16'b1011001101110000;
				18'b011000101000101111: oled_data = 16'b1010101100101111;
				18'b011000101010101111: oled_data = 16'b1010101100101111;
				18'b011000101100101111: oled_data = 16'b1011110000010010;
				18'b011000101110101111: oled_data = 16'b1101111001011001;
				18'b011000110000101111: oled_data = 16'b1110111100011011;
				18'b011000110010101111: oled_data = 16'b1110011011111010;
				18'b011000110100101111: oled_data = 16'b1110011011111010;
				18'b011000110110101111: oled_data = 16'b1110011011111010;
				18'b011000111000101111: oled_data = 16'b1110011011111010;
				18'b011000111010101111: oled_data = 16'b1110011011111010;
				18'b011000111100101111: oled_data = 16'b1110011011111010;
				18'b011000111110101111: oled_data = 16'b1110011011111010;
				18'b011001000000101111: oled_data = 16'b1110011011111010;
				18'b011001000010101111: oled_data = 16'b1110011011111010;
				18'b011001000100101111: oled_data = 16'b1110011011111010;
				18'b011001000110101111: oled_data = 16'b1110011011111010;
				18'b011001001000101111: oled_data = 16'b1110011011111010;
				18'b011001001010101111: oled_data = 16'b1110011011111010;
				18'b011001001100101111: oled_data = 16'b1110011011111010;
				18'b011001001110101111: oled_data = 16'b1110011011111010;
				18'b011001010000101111: oled_data = 16'b1110011011111010;
				18'b011001010010101111: oled_data = 16'b1110011011111010;
				18'b011001010100101111: oled_data = 16'b1110011011111010;
				18'b011001010110101111: oled_data = 16'b1110011011111010;
				18'b011001011000101111: oled_data = 16'b1110011011111010;
				18'b011001011010101111: oled_data = 16'b1110011100011010;
				18'b011001011100101111: oled_data = 16'b1110111100011010;
				18'b011001011110101111: oled_data = 16'b1101111000010111;
				18'b011001100000101111: oled_data = 16'b1011010000110001;
				18'b011001100010101111: oled_data = 16'b1100010001010001;
				18'b011001100100101111: oled_data = 16'b1101110100110101;
				18'b011001100110101111: oled_data = 16'b1101010011010011;
				18'b011001101000101111: oled_data = 16'b1101110100110101;
				18'b011001101010101111: oled_data = 16'b1101110100110101;
				18'b011001101100101111: oled_data = 16'b1101110100110101;
				18'b011001101110101111: oled_data = 16'b1101111000011000;
				18'b011001110000101111: oled_data = 16'b1110111100011010;
				18'b011001110010101111: oled_data = 16'b1101111010011000;
				18'b011001110100101111: oled_data = 16'b1110011011111010;
				18'b011001110110101111: oled_data = 16'b1110111011111010;
				18'b011001111000101111: oled_data = 16'b1110011011111010;
				18'b011001111010101111: oled_data = 16'b1110011100011010;
				18'b011001111100101111: oled_data = 16'b1110011011111001;
				18'b011001111110101111: oled_data = 16'b1010101100101100;
				18'b011010000000101111: oled_data = 16'b1011001001101010;
				18'b011010000010101111: oled_data = 16'b1100101111101111;
				18'b011010000100101111: oled_data = 16'b1011001001001001;
				18'b011010000110101111: oled_data = 16'b1011001000101001;
				18'b011010001000101111: oled_data = 16'b1011001001101001;
				18'b011010001010101111: oled_data = 16'b1011001001001001;
				18'b011010001100101111: oled_data = 16'b1011001000101000;
				18'b011010001110101111: oled_data = 16'b1011101011101100;
				18'b011010010000101111: oled_data = 16'b1100011010111011;
				18'b011010010010101111: oled_data = 16'b1011111011011100;
				18'b011010010100101111: oled_data = 16'b1011111011011011;
				18'b011010010110101111: oled_data = 16'b1011111011011011;
				18'b011010011000101111: oled_data = 16'b1011111011011011;
				18'b011010011010101111: oled_data = 16'b1100011011111100;
				18'b011010011100101111: oled_data = 16'b1011111100011100;
				18'b011010011110101111: oled_data = 16'b1011110100010100;
				18'b011010100000101111: oled_data = 16'b1010100111101000;
				18'b011010100010101111: oled_data = 16'b1010100111101000;
				18'b011010100100101111: oled_data = 16'b1010101000001000;
				18'b011010100110101111: oled_data = 16'b1010100111101000;
				18'b011000011000110000: oled_data = 16'b1010101111010001;
				18'b011000011010110000: oled_data = 16'b1101110010010101;
				18'b011000011100110000: oled_data = 16'b1101010001110100;
				18'b011000011110110000: oled_data = 16'b1100110000110011;
				18'b011000100000110000: oled_data = 16'b1101110010110101;
				18'b011000100010110000: oled_data = 16'b1011101110110001;
				18'b011000100100110000: oled_data = 16'b1010101100110000;
				18'b011000100110110000: oled_data = 16'b1011001101010000;
				18'b011000101000110000: oled_data = 16'b1010001100001111;
				18'b011000101010110000: oled_data = 16'b1011001101010000;
				18'b011000101100110000: oled_data = 16'b1010101100001111;
				18'b011000101110110000: oled_data = 16'b1011001110010000;
				18'b011000110000110000: oled_data = 16'b1101010101110110;
				18'b011000110010110000: oled_data = 16'b1110011011111010;
				18'b011000110100110000: oled_data = 16'b1110011100011010;
				18'b011000110110110000: oled_data = 16'b1110011011111010;
				18'b011000111000110000: oled_data = 16'b1110011011111010;
				18'b011000111010110000: oled_data = 16'b1110011011111010;
				18'b011000111100110000: oled_data = 16'b1110011011011001;
				18'b011000111110110000: oled_data = 16'b1110011011011001;
				18'b011001000000110000: oled_data = 16'b1110011011011001;
				18'b011001000010110000: oled_data = 16'b1110011011011001;
				18'b011001000100110000: oled_data = 16'b1110011011011010;
				18'b011001000110110000: oled_data = 16'b1110011011111010;
				18'b011001001000110000: oled_data = 16'b1110011011111010;
				18'b011001001010110000: oled_data = 16'b1110011011111010;
				18'b011001001100110000: oled_data = 16'b1110011011111010;
				18'b011001001110110000: oled_data = 16'b1110011011111010;
				18'b011001010000110000: oled_data = 16'b1110011011111010;
				18'b011001010010110000: oled_data = 16'b1110011011111010;
				18'b011001010100110000: oled_data = 16'b1110011011111010;
				18'b011001010110110000: oled_data = 16'b1110011100011010;
				18'b011001011000110000: oled_data = 16'b1110111100011010;
				18'b011001011010110000: oled_data = 16'b1110011001111000;
				18'b011001011100110000: oled_data = 16'b1100010011110011;
				18'b011001011110110000: oled_data = 16'b1011001111001111;
				18'b011001100000110000: oled_data = 16'b1011101110101111;
				18'b011001100010110000: oled_data = 16'b1101110011110100;
				18'b011001100100110000: oled_data = 16'b1101010011010100;
				18'b011001100110110000: oled_data = 16'b1101010011110100;
				18'b011001101000110000: oled_data = 16'b1101110100110101;
				18'b011001101010110000: oled_data = 16'b1101110100110101;
				18'b011001101100110000: oled_data = 16'b1101010100110101;
				18'b011001101110110000: oled_data = 16'b1100110101010101;
				18'b011001110000110000: oled_data = 16'b1101111000111000;
				18'b011001110010110000: oled_data = 16'b1110011010111001;
				18'b011001110100110000: oled_data = 16'b1110011011111010;
				18'b011001110110110000: oled_data = 16'b1110011011111010;
				18'b011001111000110000: oled_data = 16'b1110011011111010;
				18'b011001111010110000: oled_data = 16'b1110011011111010;
				18'b011001111100110000: oled_data = 16'b1110011011011001;
				18'b011001111110110000: oled_data = 16'b1011001110101110;
				18'b011010000000110000: oled_data = 16'b1011001001101010;
				18'b011010000010110000: oled_data = 16'b1100101110001110;
				18'b011010000100110000: oled_data = 16'b1011001000101001;
				18'b011010000110110000: oled_data = 16'b1011001000101001;
				18'b011010001000110000: oled_data = 16'b1100101101001101;
				18'b011010001010110000: oled_data = 16'b1011101001101010;
				18'b011010001100110000: oled_data = 16'b1011001000101000;
				18'b011010001110110000: oled_data = 16'b1011101100001100;
				18'b011010010000110000: oled_data = 16'b1100011010111011;
				18'b011010010010110000: oled_data = 16'b1011111011011100;
				18'b011010010100110000: oled_data = 16'b1011111011011100;
				18'b011010010110110000: oled_data = 16'b1011111010111011;
				18'b011010011000110000: oled_data = 16'b1011011010011010;
				18'b011010011010110000: oled_data = 16'b1011011010111011;
				18'b011010011100110000: oled_data = 16'b1011111100111100;
				18'b011010011110110000: oled_data = 16'b1011110100110101;
				18'b011010100000110000: oled_data = 16'b1010100111001000;
				18'b011010100010110000: oled_data = 16'b1001100111000111;
				18'b011010100100110000: oled_data = 16'b1001100111000111;
				18'b011010100110110000: oled_data = 16'b1001100111000111;
				18'b011000011000110001: oled_data = 16'b1001101110010000;
				18'b011000011010110001: oled_data = 16'b1101010001110100;
				18'b011000011100110001: oled_data = 16'b1101010001010100;
				18'b011000011110110001: oled_data = 16'b1100110000010011;
				18'b011000100000110001: oled_data = 16'b1101010010010101;
				18'b011000100010110001: oled_data = 16'b1011101110110001;
				18'b011000100100110001: oled_data = 16'b1010101100101111;
				18'b011000100110110001: oled_data = 16'b1010101100101111;
				18'b011000101000110001: oled_data = 16'b1010001100001110;
				18'b011000101010110001: oled_data = 16'b1010101100101111;
				18'b011000101100110001: oled_data = 16'b1010001011101110;
				18'b011000101110110001: oled_data = 16'b1010001011001110;
				18'b011000110000110001: oled_data = 16'b1001101011101110;
				18'b011000110010110001: oled_data = 16'b1010110000110001;
				18'b011000110100110001: oled_data = 16'b1101010110110110;
				18'b011000110110110001: oled_data = 16'b1110011010111001;
				18'b011000111000110001: oled_data = 16'b1110011100011010;
				18'b011000111010110001: oled_data = 16'b1110011011111010;
				18'b011000111100110001: oled_data = 16'b1110011011111010;
				18'b011000111110110001: oled_data = 16'b1110011011011010;
				18'b011001000000110001: oled_data = 16'b1110011011011001;
				18'b011001000010110001: oled_data = 16'b1110011011011001;
				18'b011001000100110001: oled_data = 16'b1110011011011010;
				18'b011001000110110001: oled_data = 16'b1110011011111010;
				18'b011001001000110001: oled_data = 16'b1110011011111010;
				18'b011001001010110001: oled_data = 16'b1110011011111010;
				18'b011001001100110001: oled_data = 16'b1110011011111010;
				18'b011001001110110001: oled_data = 16'b1110011011111010;
				18'b011001010000110001: oled_data = 16'b1110011011111010;
				18'b011001010010110001: oled_data = 16'b1110011011111010;
				18'b011001010100110001: oled_data = 16'b1110111100011010;
				18'b011001010110110001: oled_data = 16'b1110011010111001;
				18'b011001011000110001: oled_data = 16'b1100110101010100;
				18'b011001011010110001: oled_data = 16'b1011001111110000;
				18'b011001011100110001: oled_data = 16'b1011101110101111;
				18'b011001011110110001: oled_data = 16'b1011101111010000;
				18'b011001100000110001: oled_data = 16'b1100110001010010;
				18'b011001100010110001: oled_data = 16'b1101110011110100;
				18'b011001100100110001: oled_data = 16'b1101010010110011;
				18'b011001100110110001: oled_data = 16'b1101110100010101;
				18'b011001101000110001: oled_data = 16'b1101110100010101;
				18'b011001101010110001: oled_data = 16'b1101110100010101;
				18'b011001101100110001: oled_data = 16'b1101110100010101;
				18'b011001101110110001: oled_data = 16'b1101010100010100;
				18'b011001110000110001: oled_data = 16'b1100110011110100;
				18'b011001110010110001: oled_data = 16'b1101111001111001;
				18'b011001110100110001: oled_data = 16'b1110111100011010;
				18'b011001110110110001: oled_data = 16'b1110011011111010;
				18'b011001111000110001: oled_data = 16'b1110011011011010;
				18'b011001111010110001: oled_data = 16'b1110011011011001;
				18'b011001111100110001: oled_data = 16'b1101111010011000;
				18'b011001111110110001: oled_data = 16'b1011001111001110;
				18'b011010000000110001: oled_data = 16'b1011001001101001;
				18'b011010000010110001: oled_data = 16'b1100001101001101;
				18'b011010000100110001: oled_data = 16'b1011001000101001;
				18'b011010000110110001: oled_data = 16'b1011001001001001;
				18'b011010001000110001: oled_data = 16'b1100101101101101;
				18'b011010001010110001: oled_data = 16'b1011001001001001;
				18'b011010001100110001: oled_data = 16'b1011001000001000;
				18'b011010001110110001: oled_data = 16'b1011101011101011;
				18'b011010010000110001: oled_data = 16'b1100011010111011;
				18'b011010010010110001: oled_data = 16'b1011111011111100;
				18'b011010010100110001: oled_data = 16'b1011011011011011;
				18'b011010010110110001: oled_data = 16'b1001110111111001;
				18'b011010011000110001: oled_data = 16'b1001010110111000;
				18'b011010011010110001: oled_data = 16'b1010111001111010;
				18'b011010011100110001: oled_data = 16'b1011111100011100;
				18'b011010011110110001: oled_data = 16'b1011010010010010;
				18'b011010100000110001: oled_data = 16'b1010000111000111;
				18'b011010100010110001: oled_data = 16'b1010000111101000;
				18'b011010100100110001: oled_data = 16'b1010000111101000;
				18'b011010100110110001: oled_data = 16'b1010000111000111;
				18'b011000011000110010: oled_data = 16'b1000001100001101;
				18'b011000011010110010: oled_data = 16'b1101010001010100;
				18'b011000011100110010: oled_data = 16'b1101010001010100;
				18'b011000011110110010: oled_data = 16'b1100001111110010;
				18'b011000100000110010: oled_data = 16'b1100110001010100;
				18'b011000100010110010: oled_data = 16'b1011101110010001;
				18'b011000100100110010: oled_data = 16'b1010101100101111;
				18'b011000100110110010: oled_data = 16'b1010001011101110;
				18'b011000101000110010: oled_data = 16'b1010001011101110;
				18'b011000101010110010: oled_data = 16'b1010101100001111;
				18'b011000101100110010: oled_data = 16'b1001101011001110;
				18'b011000101110110010: oled_data = 16'b1001101011001110;
				18'b011000110000110010: oled_data = 16'b1010001011101110;
				18'b011000110010110010: oled_data = 16'b1010101100101111;
				18'b011000110100110010: oled_data = 16'b1010101101001111;
				18'b011000110110110010: oled_data = 16'b1011001111110000;
				18'b011000111000110010: oled_data = 16'b1011110011110011;
				18'b011000111010110010: oled_data = 16'b1101010110110110;
				18'b011000111100110010: oled_data = 16'b1101111001111000;
				18'b011000111110110010: oled_data = 16'b1110111011011010;
				18'b011001000000110010: oled_data = 16'b1110111011111010;
				18'b011001000010110010: oled_data = 16'b1110011011111010;
				18'b011001000100110010: oled_data = 16'b1110011011111010;
				18'b011001000110110010: oled_data = 16'b1110011011111010;
				18'b011001001000110010: oled_data = 16'b1110011011011001;
				18'b011001001010110010: oled_data = 16'b1101111010111001;
				18'b011001001100110010: oled_data = 16'b1101111011011001;
				18'b011001001110110010: oled_data = 16'b1110011011111010;
				18'b011001010000110010: oled_data = 16'b1101111010111001;
				18'b011001010010110010: oled_data = 16'b1101010111010110;
				18'b011001010100110010: oled_data = 16'b1100010011110011;
				18'b011001010110110010: oled_data = 16'b1011001111110000;
				18'b011001011000110010: oled_data = 16'b1011001110001111;
				18'b011001011010110010: oled_data = 16'b1011101110110000;
				18'b011001011100110010: oled_data = 16'b1011101111010000;
				18'b011001011110110010: oled_data = 16'b1100110001010010;
				18'b011001100000110010: oled_data = 16'b1101010010110011;
				18'b011001100010110010: oled_data = 16'b1100110010010011;
				18'b011001100100110010: oled_data = 16'b1101010011110100;
				18'b011001100110110010: oled_data = 16'b1101110100010101;
				18'b011001101000110010: oled_data = 16'b1101110100010101;
				18'b011001101010110010: oled_data = 16'b1101110100010101;
				18'b011001101100110010: oled_data = 16'b1101110100010101;
				18'b011001101110110010: oled_data = 16'b1101010011110100;
				18'b011001110000110010: oled_data = 16'b1101010011110100;
				18'b011001110010110010: oled_data = 16'b1100110011110100;
				18'b011001110100110010: oled_data = 16'b1100110110010101;
				18'b011001110110110010: oled_data = 16'b1101111010111001;
				18'b011001111000110010: oled_data = 16'b1110011011111010;
				18'b011001111010110010: oled_data = 16'b1110011011011010;
				18'b011001111100110010: oled_data = 16'b1110011011011010;
				18'b011001111110110010: oled_data = 16'b1011001111001110;
				18'b011010000000110010: oled_data = 16'b1011001001001001;
				18'b011010000010110010: oled_data = 16'b1100001100101100;
				18'b011010000100110010: oled_data = 16'b1011001000101001;
				18'b011010000110110010: oled_data = 16'b1011001001001001;
				18'b011010001000110010: oled_data = 16'b1011101010101010;
				18'b011010001010110010: oled_data = 16'b1011001000101000;
				18'b011010001100110010: oled_data = 16'b1011001000001000;
				18'b011010001110110010: oled_data = 16'b1011001001101010;
				18'b011010010000110010: oled_data = 16'b1100011001011001;
				18'b011010010010110010: oled_data = 16'b1011111011111100;
				18'b011010010100110010: oled_data = 16'b1010011000111001;
				18'b011010010110110010: oled_data = 16'b1001010110110111;
				18'b011010011000110010: oled_data = 16'b1001010110111000;
				18'b011010011010110010: oled_data = 16'b1001110111111000;
				18'b011010011100110010: oled_data = 16'b1010111010011010;
				18'b011010011110110010: oled_data = 16'b1010101110101111;
				18'b011010100000110010: oled_data = 16'b1010000110100111;
				18'b011010100010110010: oled_data = 16'b1010000111000111;
				18'b011010100100110010: oled_data = 16'b1010000111000111;
				18'b011010100110110010: oled_data = 16'b1010000111000111;
				18'b011000011000110011: oled_data = 16'b0110001001101010;
				18'b011000011010110011: oled_data = 16'b1100110000110011;
				18'b011000011100110011: oled_data = 16'b1100110000110011;
				18'b011000011110110011: oled_data = 16'b1100001111110011;
				18'b011000100000110011: oled_data = 16'b1100001111110011;
				18'b011000100010110011: oled_data = 16'b1011101111010001;
				18'b011000100100110011: oled_data = 16'b1010101100101111;
				18'b011000100110110011: oled_data = 16'b1001101010101101;
				18'b011000101000110011: oled_data = 16'b1010001011101111;
				18'b011000101010110011: oled_data = 16'b1010001011101110;
				18'b011000101100110011: oled_data = 16'b1001101010101101;
				18'b011000101110110011: oled_data = 16'b1001101010001101;
				18'b011000110000110011: oled_data = 16'b1010001011101110;
				18'b011000110010110011: oled_data = 16'b1010101100101111;
				18'b011000110100110011: oled_data = 16'b1010101100101110;
				18'b011000110110110011: oled_data = 16'b1010101100101110;
				18'b011000111000110011: oled_data = 16'b1010001100101110;
				18'b011000111010110011: oled_data = 16'b1010001100101110;
				18'b011000111100110011: oled_data = 16'b1010101110001111;
				18'b011000111110110011: oled_data = 16'b1011010000110001;
				18'b011001000000110011: oled_data = 16'b1100010011110100;
				18'b011001000010110011: oled_data = 16'b1100010101110101;
				18'b011001000100110011: oled_data = 16'b1101010111010110;
				18'b011001000110110011: oled_data = 16'b1100110111010110;
				18'b011001001000110011: oled_data = 16'b1101011000110111;
				18'b011001001010110011: oled_data = 16'b1101011001111000;
				18'b011001001100110011: oled_data = 16'b1101011001010111;
				18'b011001001110110011: oled_data = 16'b1011010011010010;
				18'b011001010000110011: oled_data = 16'b1010101110101111;
				18'b011001010010110011: oled_data = 16'b1011001110001111;
				18'b011001010100110011: oled_data = 16'b1011001101101111;
				18'b011001010110110011: oled_data = 16'b1011001101101111;
				18'b011001011000110011: oled_data = 16'b1011001110001111;
				18'b011001011010110011: oled_data = 16'b1011001110101111;
				18'b011001011100110011: oled_data = 16'b1100010000110001;
				18'b011001011110110011: oled_data = 16'b1101010010110011;
				18'b011001100000110011: oled_data = 16'b1100010000110001;
				18'b011001100010110011: oled_data = 16'b1101010011010100;
				18'b011001100100110011: oled_data = 16'b1101110011110100;
				18'b011001100110110011: oled_data = 16'b1101010011110100;
				18'b011001101000110011: oled_data = 16'b1101110011110101;
				18'b011001101010110011: oled_data = 16'b1101010011110100;
				18'b011001101100110011: oled_data = 16'b1101010011110100;
				18'b011001101110110011: oled_data = 16'b1101010011110100;
				18'b011001110000110011: oled_data = 16'b1101010011010100;
				18'b011001110010110011: oled_data = 16'b1101010011010100;
				18'b011001110100110011: oled_data = 16'b0110001000001000;
				18'b011001110110110011: oled_data = 16'b0100101000100111;
				18'b011001111000110011: oled_data = 16'b1011010101110100;
				18'b011001111010110011: oled_data = 16'b1101111010111010;
				18'b011001111100110011: oled_data = 16'b1010010011010001;
				18'b011001111110110011: oled_data = 16'b1000101001001000;
				18'b011010000000110011: oled_data = 16'b1011101001101010;
				18'b011010000010110011: oled_data = 16'b1011101100001100;
				18'b011010000100110011: oled_data = 16'b1011001000001000;
				18'b011010000110110011: oled_data = 16'b1011001000001000;
				18'b011010001000110011: oled_data = 16'b1011001000001000;
				18'b011010001010110011: oled_data = 16'b1011001000001000;
				18'b011010001100110011: oled_data = 16'b1010101000001000;
				18'b011010001110110011: oled_data = 16'b1011001000001000;
				18'b011010010000110011: oled_data = 16'b1011110100010100;
				18'b011010010010110011: oled_data = 16'b1011011011111011;
				18'b011010010100110011: oled_data = 16'b1001010111010111;
				18'b011010010110110011: oled_data = 16'b1000110110010110;
				18'b011010011000110011: oled_data = 16'b1000110110010110;
				18'b011010011010110011: oled_data = 16'b1000110110010111;
				18'b011010011100110011: oled_data = 16'b1010010111010111;
				18'b011010011110110011: oled_data = 16'b1010001001101010;
				18'b011010100000110011: oled_data = 16'b1010000111000111;
				18'b011010100010110011: oled_data = 16'b1010000111000111;
				18'b011010100100110011: oled_data = 16'b1001100111000111;
				18'b011010100110110011: oled_data = 16'b1001100111000111;
				18'b011000011000110100: oled_data = 16'b0100000111001000;
				18'b011000011010110100: oled_data = 16'b1011001111010001;
				18'b011000011100110100: oled_data = 16'b1100110000010011;
				18'b011000011110110100: oled_data = 16'b1100110000010011;
				18'b011000100000110100: oled_data = 16'b1011101110110001;
				18'b011000100010110100: oled_data = 16'b1011101111010010;
				18'b011000100100110100: oled_data = 16'b1100001111010010;
				18'b011000100110110100: oled_data = 16'b1010001011101110;
				18'b011000101000110100: oled_data = 16'b1001101010101110;
				18'b011000101010110100: oled_data = 16'b1010001011101110;
				18'b011000101100110100: oled_data = 16'b1001001010001101;
				18'b011000101110110100: oled_data = 16'b1001001001101100;
				18'b011000110000110100: oled_data = 16'b1010101100101111;
				18'b011000110010110100: oled_data = 16'b1010101101001111;
				18'b011000110100110100: oled_data = 16'b1010001100001110;
				18'b011000110110110100: oled_data = 16'b1010101101001110;
				18'b011000111000110100: oled_data = 16'b1010101101101111;
				18'b011000111010110100: oled_data = 16'b1011001110110000;
				18'b011000111100110100: oled_data = 16'b1011001110110000;
				18'b011000111110110100: oled_data = 16'b1011001110010000;
				18'b011001000000110100: oled_data = 16'b1010101101101111;
				18'b011001000010110100: oled_data = 16'b1010001101001110;
				18'b011001000100110100: oled_data = 16'b1010001100101110;
				18'b011001000110110100: oled_data = 16'b1011010001110010;
				18'b011001001000110100: oled_data = 16'b1101111001111000;
				18'b011001001010110100: oled_data = 16'b1101111010111001;
				18'b011001001100110100: oled_data = 16'b1101111010111001;
				18'b011001001110110100: oled_data = 16'b1101011000010111;
				18'b011001010000110100: oled_data = 16'b1011010001010001;
				18'b011001010010110100: oled_data = 16'b1011001101101111;
				18'b011001010100110100: oled_data = 16'b1011001101101110;
				18'b011001010110110100: oled_data = 16'b1010101100101101;
				18'b011001011000110100: oled_data = 16'b1011001110101111;
				18'b011001011010110100: oled_data = 16'b1100010000110001;
				18'b011001011100110100: oled_data = 16'b1100110001010010;
				18'b011001011110110100: oled_data = 16'b1101010010010011;
				18'b011001100000110100: oled_data = 16'b1100110001010010;
				18'b011001100010110100: oled_data = 16'b1101010010110100;
				18'b011001100100110100: oled_data = 16'b1101010011010100;
				18'b011001100110110100: oled_data = 16'b1101010011010100;
				18'b011001101000110100: oled_data = 16'b1101010011010100;
				18'b011001101010110100: oled_data = 16'b1101010011010100;
				18'b011001101100110100: oled_data = 16'b1101010011010100;
				18'b011001101110110100: oled_data = 16'b1101010011010100;
				18'b011001110000110100: oled_data = 16'b1101010011010100;
				18'b011001110010110100: oled_data = 16'b1011110001010010;
				18'b011001110100110100: oled_data = 16'b0011000011100011;
				18'b011001110110110100: oled_data = 16'b0001000010000001;
				18'b011001111000110100: oled_data = 16'b0010000100000011;
				18'b011001111010110100: oled_data = 16'b0100000111100111;
				18'b011001111100110100: oled_data = 16'b0010000011000010;
				18'b011001111110110100: oled_data = 16'b0111000110000101;
				18'b011010000000110100: oled_data = 16'b1011101001001010;
				18'b011010000010110100: oled_data = 16'b1011001011001011;
				18'b011010000100110100: oled_data = 16'b1010101000001000;
				18'b011010000110110100: oled_data = 16'b1010101000001000;
				18'b011010001000110100: oled_data = 16'b1010101000001000;
				18'b011010001010110100: oled_data = 16'b1010101000001000;
				18'b011010001100110100: oled_data = 16'b1010101000001000;
				18'b011010001110110100: oled_data = 16'b1010100111101000;
				18'b011010010000110100: oled_data = 16'b1001101001001010;
				18'b011010010010110100: oled_data = 16'b1011111000011000;
				18'b011010010100110100: oled_data = 16'b1001111000111000;
				18'b011010010110110100: oled_data = 16'b1000110110010110;
				18'b011010011000110100: oled_data = 16'b1000110110010111;
				18'b011010011010110100: oled_data = 16'b1001010110110111;
				18'b011010011100110100: oled_data = 16'b1010001110101111;
				18'b011010011110110100: oled_data = 16'b1001100110100111;
				18'b011010100000110100: oled_data = 16'b1010000111000111;
				18'b011010100010110100: oled_data = 16'b1001100110100111;
				18'b011010100100110100: oled_data = 16'b1001100110100111;
				18'b011010100110110100: oled_data = 16'b1001100110100111;
				18'b011000011000110101: oled_data = 16'b0011000101100110;
				18'b011000011010110101: oled_data = 16'b1000101011001101;
				18'b011000011100110101: oled_data = 16'b1100110000010011;
				18'b011000011110110101: oled_data = 16'b1100001111110010;
				18'b011000100000110101: oled_data = 16'b1011101110110001;
				18'b011000100010110101: oled_data = 16'b1011101110010001;
				18'b011000100100110101: oled_data = 16'b1100001111110010;
				18'b011000100110110101: oled_data = 16'b1100001111010010;
				18'b011000101000110101: oled_data = 16'b1010001011001110;
				18'b011000101010110101: oled_data = 16'b1001101010101101;
				18'b011000101100110101: oled_data = 16'b1000101001001100;
				18'b011000101110110101: oled_data = 16'b1001101010001100;
				18'b011000110000110101: oled_data = 16'b1010101100101110;
				18'b011000110010110101: oled_data = 16'b1010101100101110;
				18'b011000110100110101: oled_data = 16'b1011001110110000;
				18'b011000110110110101: oled_data = 16'b1100010000110010;
				18'b011000111000110101: oled_data = 16'b1100110001110011;
				18'b011000111010110101: oled_data = 16'b1100110010010011;
				18'b011000111100110101: oled_data = 16'b1100110010010011;
				18'b011000111110110101: oled_data = 16'b1100110001110011;
				18'b011001000000110101: oled_data = 16'b1011110000010001;
				18'b011001000010110101: oled_data = 16'b1010101110001111;
				18'b011001000100110101: oled_data = 16'b1010110000110001;
				18'b011001000110110101: oled_data = 16'b1101111001111001;
				18'b011001001000110101: oled_data = 16'b1101111010011001;
				18'b011001001010110101: oled_data = 16'b1101111010011000;
				18'b011001001100110101: oled_data = 16'b1101111010011000;
				18'b011001001110110101: oled_data = 16'b1101111010011001;
				18'b011001010000110101: oled_data = 16'b1101111001011000;
				18'b011001010010110101: oled_data = 16'b1011110000010001;
				18'b011001010100110101: oled_data = 16'b1100110000010001;
				18'b011001010110110101: oled_data = 16'b1100110001110010;
				18'b011001011000110101: oled_data = 16'b1101010010010011;
				18'b011001011010110101: oled_data = 16'b1101010010110011;
				18'b011001011100110101: oled_data = 16'b1101010010110011;
				18'b011001011110110101: oled_data = 16'b1101010010110011;
				18'b011001100000110101: oled_data = 16'b1100010001010010;
				18'b011001100010110101: oled_data = 16'b1100110010010011;
				18'b011001100100110101: oled_data = 16'b1101010010110100;
				18'b011001100110110101: oled_data = 16'b1101010010110100;
				18'b011001101000110101: oled_data = 16'b1101010010110100;
				18'b011001101010110101: oled_data = 16'b1100110010110011;
				18'b011001101100110101: oled_data = 16'b1100110010110011;
				18'b011001101110110101: oled_data = 16'b1100110010110011;
				18'b011001110000110101: oled_data = 16'b1101010011010100;
				18'b011001110010110101: oled_data = 16'b1001001101001110;
				18'b011001110100110101: oled_data = 16'b0001100001100001;
				18'b011001110110110101: oled_data = 16'b0001100010000001;
				18'b011001111000110101: oled_data = 16'b0010000010100010;
				18'b011001111010110101: oled_data = 16'b0010100011000010;
				18'b011001111100110101: oled_data = 16'b0100000100100100;
				18'b011001111110110101: oled_data = 16'b0111100111000110;
				18'b011010000000110101: oled_data = 16'b1011001000001001;
				18'b011010000010110101: oled_data = 16'b1011001010001010;
				18'b011010000100110101: oled_data = 16'b1010101000001000;
				18'b011010000110110101: oled_data = 16'b1010101000001000;
				18'b011010001000110101: oled_data = 16'b1010101000001000;
				18'b011010001010110101: oled_data = 16'b1010101000001000;
				18'b011010001100110101: oled_data = 16'b1010100111101000;
				18'b011010001110110101: oled_data = 16'b1010000111101000;
				18'b011010010000110101: oled_data = 16'b1000100101000110;
				18'b011010010010110101: oled_data = 16'b1010101011001100;
				18'b011010010100110101: oled_data = 16'b1011010011010011;
				18'b011010010110110101: oled_data = 16'b1010010011110011;
				18'b011010011000110101: oled_data = 16'b1010010001010010;
				18'b011010011010110101: oled_data = 16'b1010001101001110;
				18'b011010011100110101: oled_data = 16'b1001100111101000;
				18'b011010011110110101: oled_data = 16'b1010000111000111;
				18'b011010100000110101: oled_data = 16'b1001100111000111;
				18'b011010100010110101: oled_data = 16'b1001100110100111;
				18'b011010100100110101: oled_data = 16'b1001100110100111;
				18'b011010100110110101: oled_data = 16'b1001100110100111;
				18'b011000011000110110: oled_data = 16'b0010100101100110;
				18'b011000011010110110: oled_data = 16'b0110101001001011;
				18'b011000011100110110: oled_data = 16'b1100001111010010;
				18'b011000011110110110: oled_data = 16'b1100001111010010;
				18'b011000100000110110: oled_data = 16'b1011101110110001;
				18'b011000100010110110: oled_data = 16'b1011001101010000;
				18'b011000100100110110: oled_data = 16'b1011101110110001;
				18'b011000100110110110: oled_data = 16'b1100110000010011;
				18'b011000101000110110: oled_data = 16'b1100001111010010;
				18'b011000101010110110: oled_data = 16'b1010101101010000;
				18'b011000101100110110: oled_data = 16'b1000101000101011;
				18'b011000101110110110: oled_data = 16'b1001001010001100;
				18'b011000110000110110: oled_data = 16'b1011001101001111;
				18'b011000110010110110: oled_data = 16'b1100010000010010;
				18'b011000110100110110: oled_data = 16'b1100110001010010;
				18'b011000110110110110: oled_data = 16'b1100010001010011;
				18'b011000111000110110: oled_data = 16'b1100110001110011;
				18'b011000111010110110: oled_data = 16'b1100110001110011;
				18'b011000111100110110: oled_data = 16'b1100110001010011;
				18'b011000111110110110: oled_data = 16'b1100010001010010;
				18'b011001000000110110: oled_data = 16'b1100010000110001;
				18'b011001000010110110: oled_data = 16'b1011010000110001;
				18'b011001000100110110: oled_data = 16'b1100111000010111;
				18'b011001000110110110: oled_data = 16'b1101011001111000;
				18'b011001001000110110: oled_data = 16'b1101011001111000;
				18'b011001001010110110: oled_data = 16'b1101011001011000;
				18'b011001001100110110: oled_data = 16'b1101011001010111;
				18'b011001001110110110: oled_data = 16'b1101011001011000;
				18'b011001010000110110: oled_data = 16'b1101011001111000;
				18'b011001010010110110: oled_data = 16'b1100010100110100;
				18'b011001010100110110: oled_data = 16'b1100110001110010;
				18'b011001010110110110: oled_data = 16'b1100110001110010;
				18'b011001011000110110: oled_data = 16'b1100110010010010;
				18'b011001011010110110: oled_data = 16'b1100110010010011;
				18'b011001011100110110: oled_data = 16'b1100110010010011;
				18'b011001011110110110: oled_data = 16'b1101010010010011;
				18'b011001100000110110: oled_data = 16'b1100010000110010;
				18'b011001100010110110: oled_data = 16'b1100110001110011;
				18'b011001100100110110: oled_data = 16'b1100110010010100;
				18'b011001100110110110: oled_data = 16'b1100110010010100;
				18'b011001101000110110: oled_data = 16'b1100110010010011;
				18'b011001101010110110: oled_data = 16'b1100110010010011;
				18'b011001101100110110: oled_data = 16'b1100110010010011;
				18'b011001101110110110: oled_data = 16'b1100110010010011;
				18'b011001110000110110: oled_data = 16'b1100110010010011;
				18'b011001110010110110: oled_data = 16'b0101100110100111;
				18'b011001110100110110: oled_data = 16'b0010000001100001;
				18'b011001110110110110: oled_data = 16'b0010100010100010;
				18'b011001111000110110: oled_data = 16'b0011100100000011;
				18'b011001111010110110: oled_data = 16'b0101100111000101;
				18'b011001111100110110: oled_data = 16'b0111101001101000;
				18'b011001111110110110: oled_data = 16'b1001001000100111;
				18'b011010000000110110: oled_data = 16'b1011001000001000;
				18'b011010000010110110: oled_data = 16'b1010101001101001;
				18'b011010000100110110: oled_data = 16'b1010100111101000;
				18'b011010000110110110: oled_data = 16'b1010100111101000;
				18'b011010001000110110: oled_data = 16'b1010100111101000;
				18'b011010001010110110: oled_data = 16'b1010100111101000;
				18'b011010001100110110: oled_data = 16'b1010000111100111;
				18'b011010001110110110: oled_data = 16'b1001100111000111;
				18'b011010010000110110: oled_data = 16'b1000100110000110;
				18'b011010010010110110: oled_data = 16'b1010000111000111;
				18'b011010010100110110: oled_data = 16'b1010000111001000;
				18'b011010010110110110: oled_data = 16'b1010000111101000;
				18'b011010011000110110: oled_data = 16'b1001100110100111;
				18'b011010011010110110: oled_data = 16'b1010000110100111;
				18'b011010011100110110: oled_data = 16'b1001100111000111;
				18'b011010011110110110: oled_data = 16'b1001100110100111;
				18'b011010100000110110: oled_data = 16'b1001100110100111;
				18'b011010100010110110: oled_data = 16'b1001100110100110;
				18'b011010100100110110: oled_data = 16'b1001000110000110;
				18'b011010100110110110: oled_data = 16'b1001000110000110;
				18'b011000011000110111: oled_data = 16'b0010100100100101;
				18'b011000011010110111: oled_data = 16'b0111101001001011;
				18'b011000011100110111: oled_data = 16'b1011101101010000;
				18'b011000011110110111: oled_data = 16'b1100001110110001;
				18'b011000100000110111: oled_data = 16'b1100001110110001;
				18'b011000100010110111: oled_data = 16'b1011101101010000;
				18'b011000100100110111: oled_data = 16'b1011001101110000;
				18'b011000100110110111: oled_data = 16'b1100001111010010;
				18'b011000101000110111: oled_data = 16'b1100001111010010;
				18'b011000101010110111: oled_data = 16'b1100001111010010;
				18'b011000101100110111: oled_data = 16'b1011001101110000;
				18'b011000101110110111: oled_data = 16'b1010001011101110;
				18'b011000110000110111: oled_data = 16'b1011101110010001;
				18'b011000110010110111: oled_data = 16'b1100001111010010;
				18'b011000110100110111: oled_data = 16'b1100010000010010;
				18'b011000110110110111: oled_data = 16'b1100110000110010;
				18'b011000111000110111: oled_data = 16'b1100010000110010;
				18'b011000111010110111: oled_data = 16'b1100010000110010;
				18'b011000111100110111: oled_data = 16'b1100001111110010;
				18'b011000111110110111: oled_data = 16'b1100001111110010;
				18'b011001000000110111: oled_data = 16'b1011101111010001;
				18'b011001000010110111: oled_data = 16'b1011010011110011;
				18'b011001000100110111: oled_data = 16'b1101011001111000;
				18'b011001000110110111: oled_data = 16'b1100111001010111;
				18'b011001001000110111: oled_data = 16'b1100111001010111;
				18'b011001001010110111: oled_data = 16'b1100111001010111;
				18'b011001001100110111: oled_data = 16'b1100010111110110;
				18'b011001001110110111: oled_data = 16'b1100010111010110;
				18'b011001010000110111: oled_data = 16'b1100111000110111;
				18'b011001010010110111: oled_data = 16'b1100110101110101;
				18'b011001010100110111: oled_data = 16'b1100010001010010;
				18'b011001010110110111: oled_data = 16'b1100110001110010;
				18'b011001011000110111: oled_data = 16'b1100110001110010;
				18'b011001011010110111: oled_data = 16'b1100110001110010;
				18'b011001011100110111: oled_data = 16'b1100110001110010;
				18'b011001011110110111: oled_data = 16'b1100110001110010;
				18'b011001100000110111: oled_data = 16'b1100010000010001;
				18'b011001100010110111: oled_data = 16'b1100010001010010;
				18'b011001100100110111: oled_data = 16'b1100110001110010;
				18'b011001100110110111: oled_data = 16'b1100110001110010;
				18'b011001101000110111: oled_data = 16'b1100110001110010;
				18'b011001101010110111: oled_data = 16'b1100110001110010;
				18'b011001101100110111: oled_data = 16'b1100110001110011;
				18'b011001101110110111: oled_data = 16'b1100110001110011;
				18'b011001110000110111: oled_data = 16'b1011001111110001;
				18'b011001110010110111: oled_data = 16'b0011000010100011;
				18'b011001110100110111: oled_data = 16'b0011000011100011;
				18'b011001110110110111: oled_data = 16'b0101000101100101;
				18'b011001111000110111: oled_data = 16'b0111001001000111;
				18'b011001111010110111: oled_data = 16'b1000001010100111;
				18'b011001111100110111: oled_data = 16'b1000001010100111;
				18'b011001111110110111: oled_data = 16'b1001101001001000;
				18'b011010000000110111: oled_data = 16'b1010100111101000;
				18'b011010000010110111: oled_data = 16'b1010001000101000;
				18'b011010000100110111: oled_data = 16'b1010100111101000;
				18'b011010000110110111: oled_data = 16'b1010100111100111;
				18'b011010001000110111: oled_data = 16'b1010000111100111;
				18'b011010001010110111: oled_data = 16'b1010000111100111;
				18'b011010001100110111: oled_data = 16'b1010000111100111;
				18'b011010001110110111: oled_data = 16'b1001100110100111;
				18'b011010010000110111: oled_data = 16'b1000100110000111;
				18'b011010010010110111: oled_data = 16'b1010000111001000;
				18'b011010010100110111: oled_data = 16'b1010000111000111;
				18'b011010010110110111: oled_data = 16'b1001100110100111;
				18'b011010011000110111: oled_data = 16'b1001000110100110;
				18'b011010011010110111: oled_data = 16'b1001100110100111;
				18'b011010011100110111: oled_data = 16'b1001100110100111;
				18'b011010011110110111: oled_data = 16'b1001100110100111;
				18'b011010100000110111: oled_data = 16'b1001100110000110;
				18'b011010100010110111: oled_data = 16'b1001000110000110;
				18'b011010100100110111: oled_data = 16'b1001000110000110;
				18'b011010100110110111: oled_data = 16'b1001000110000110;
				default: oled_data = 16'b0;
			endcase
		end
	end

	always @ (posedge clock) begin
		COUNT <= (COUNT >= ((100000000) / (frame_rate * 2)) - 1) ? 32'b0 : COUNT + 1;
		slow_clk <= (COUNT >= ((100000000) / (frame_rate * 2)) - 1) ? ~slow_clk : slow_clk;
	end

	always @ (posedge slow_clk) begin
		frame_no <= (frame_no >= 4'd6) ? 4'd1 : frame_no + 1;
	end

endmodule