`timescale 1ns / 1ps

module test (
	input clock, btnL, btnR, btnU, btnD,
	input [6:0] x, y,
	output reg [15:0] oled_data = 0,
	input [3:0] machine_state,
	output reg [3:0] menu_state = 4'd1
	);

	wire sel1 = (x >= 24 && x <= 39 && y >= 24 && y <= 39);
	wire sel2 = (x >= 40 && x <= 55 && y >= 24 && y <= 39);
	wire sel3 = (x >= 56 && x <= 71 && y >= 24 && y <= 39);
	wire sel4 = (x >= 32 && x <= 47 && y >= 41 && y <= 56);
	wire sel5 = (x >= 48 && x <= 63 && y >= 41 && y <= 56);
	
	wire sel6 = (x >= 32 && x <= 47 && y >= 24 && y <= 39);
	wire sel7 = (x >= 48 && x <= 63 && y >= 24 && y <= 39);
	wire sel8 = (x >= 32 && x <= 47 && y >= 24 && y <= 39);
	wire sel9 = (x >= 48 && x <= 63 && y >= 41 && y <= 56);

	// Edge Detection
	reg [31:0] release_count = 0;
	reg [1:0] btnL_state = 0;
	reg [1:0] btnR_state = 0;
	reg [1:0] btnU_state = 0;
	reg [1:0] btnD_state = 0;

	always @ (posedge clock) begin
		if (machine_state == 4'd0) begin
			// Left button
			if (btnL && btnL_state == 2'b0)
				btnL_state = 2'b01;
			if (btnL_state == 2'b01) begin
				if (!btnL) begin
					release_count = release_count + 1;
					if (release_count == 31'd6_250_000)
						btnL_state = 2'b10;
				end
				else
					release_count = 0;
			end
			if (btnL_state == 2'b10) begin
				btnL_state = 2'b0;
				menu_state <= (menu_state == 4'd1) ? 4'd1 : (menu_state - 4'd1);
			end

			// Right button
			if (btnR && btnR_state == 2'b0)
				btnR_state = 2'b01;
			if (btnR_state == 2'b01) begin
				if (!btnR) begin
					release_count = release_count + 1;
					if (release_count == 31'd6_250_000)
						btnR_state = 2'b10;
				end
				else
					release_count = 0;
			end
			if (btnR_state == 2'b10) begin
				btnR_state = 2'b0;
				menu_state <= (menu_state == 4'd9) ? 4'd9 : (menu_state + 4'd1);
			end

			// Up button
			if (btnU && btnU_state == 2'b0)
				btnU_state = 2'b01;
			if (btnU_state == 2'b01) begin
				if (!btnU) begin
					release_count = release_count + 1;
					if (release_count == 31'd6_250_000)
						btnU_state = 2'b10;
				end
				else
					release_count = 0;
			end
			if (btnU_state == 2'b10) begin
				btnU_state = 2'b0;
				menu_state <= (menu_state > 4'd5) ? 4'd5 : 4'd1;
			end

			// Down button
			if (btnD && btnD_state == 2'b0)
				btnD_state = 2'b01;
			if (btnD_state == 2'b01) begin
				if (!btnD) begin
					release_count = release_count + 1;
					if (release_count == 31'd6_250_000)
						btnD_state = 2'b10;
				end
				else
					release_count = 0;
			end
			if (btnD_state == 2'b10) begin
				btnD_state = 2'b0;
				menu_state <= (menu_state < 4'd6) ? 4'd6 : 4'd9;
			end
		end
	end

	always @ (*) begin
		if (machine_state == 4'b0) begin
			case ({x, y})
				14'b00000000000000: oled_data = 16'b1111111111111111;
				14'b00000010000000: oled_data = 16'b1111111111111111;
				14'b00000100000000: oled_data = 16'b1111111111111111;
				14'b00000110000000: oled_data = 16'b1111111111111111;
				14'b00001000000000: oled_data = 16'b1111111111111111;
				14'b00001010000000: oled_data = 16'b1111111111111111;
				14'b00001100000000: oled_data = 16'b1111111111111111;
				14'b00001110000000: oled_data = 16'b1111111111111111;
				14'b00010000000000: oled_data = 16'b1111111111111111;
				14'b00010010000000: oled_data = 16'b1111111111111111;
				14'b00010100000000: oled_data = 16'b1111111111111111;
				14'b00010110000000: oled_data = 16'b1111111111111111;
				14'b00011000000000: oled_data = 16'b1111111111111111;
				14'b00011010000000: oled_data = 16'b1111111111111111;
				14'b00011100000000: oled_data = 16'b1111111111111111;
				14'b00011110000000: oled_data = 16'b1111111111111111;
				14'b00100000000000: oled_data = 16'b1111111111111111;
				14'b00100010000000: oled_data = 16'b1111111111111111;
				14'b00100100000000: oled_data = 16'b1111111111111111;
				14'b00100110000000: oled_data = 16'b1111111111111111;
				14'b00101000000000: oled_data = 16'b1111111111111111;
				14'b00101010000000: oled_data = 16'b1111111111111111;
				14'b00101100000000: oled_data = 16'b1111111111111111;
				14'b00101110000000: oled_data = 16'b1111111111111111;
				14'b00110000000000: oled_data = 16'b1111111111111111;
				14'b00110010000000: oled_data = 16'b1111111111111111;
				14'b00110100000000: oled_data = 16'b1111111111111111;
				14'b00110110000000: oled_data = 16'b1111111111111111;
				14'b00111000000000: oled_data = 16'b1111111111111111;
				14'b00111010000000: oled_data = 16'b1111111111111111;
				14'b00111100000000: oled_data = 16'b1111111111111111;
				14'b00111110000000: oled_data = 16'b1111111111111111;
				14'b01000000000000: oled_data = 16'b1111111111111111;
				14'b01000010000000: oled_data = 16'b1111111111111111;
				14'b01000100000000: oled_data = 16'b1111111111111111;
				14'b01000110000000: oled_data = 16'b1111111111111111;
				14'b01001000000000: oled_data = 16'b1111111111111111;
				14'b01001010000000: oled_data = 16'b1111111111111111;
				14'b01001100000000: oled_data = 16'b1111111111111111;
				14'b01001110000000: oled_data = 16'b1111111111111111;
				14'b01010000000000: oled_data = 16'b1111111111111111;
				14'b01010010000000: oled_data = 16'b1111111111111111;
				14'b01010100000000: oled_data = 16'b1111111111111111;
				14'b01010110000000: oled_data = 16'b1111111111111111;
				14'b01011000000000: oled_data = 16'b1111111111111111;
				14'b01011010000000: oled_data = 16'b1111111111111111;
				14'b01011100000000: oled_data = 16'b1111111111111111;
				14'b01011110000000: oled_data = 16'b1111111111111111;
				14'b01100000000000: oled_data = 16'b1111111111111111;
				14'b01100010000000: oled_data = 16'b1111111111111111;
				14'b01100100000000: oled_data = 16'b1111111111111111;
				14'b01100110000000: oled_data = 16'b1111111111111111;
				14'b01101000000000: oled_data = 16'b1111111111111111;
				14'b01101010000000: oled_data = 16'b1111111111111111;
				14'b01101100000000: oled_data = 16'b1111111111111111;
				14'b01101110000000: oled_data = 16'b1111111111111111;
				14'b01110000000000: oled_data = 16'b1111111111111111;
				14'b01110010000000: oled_data = 16'b1111111111111111;
				14'b01110100000000: oled_data = 16'b1111111111111111;
				14'b01110110000000: oled_data = 16'b1111111111111111;
				14'b01111000000000: oled_data = 16'b1111111111111111;
				14'b01111010000000: oled_data = 16'b1111111111111111;
				14'b01111100000000: oled_data = 16'b1111111111111111;
				14'b01111110000000: oled_data = 16'b1111111111111111;
				14'b10000000000000: oled_data = 16'b1111111111111111;
				14'b10000010000000: oled_data = 16'b1111111111111111;
				14'b10000100000000: oled_data = 16'b1111111111111111;
				14'b10000110000000: oled_data = 16'b1111111111111111;
				14'b10001000000000: oled_data = 16'b1111111111111111;
				14'b10001010000000: oled_data = 16'b1111111111111111;
				14'b10001100000000: oled_data = 16'b1111111111111111;
				14'b10001110000000: oled_data = 16'b1111111111111111;
				14'b10010000000000: oled_data = 16'b1111111111111111;
				14'b10010010000000: oled_data = 16'b1111111111111111;
				14'b10010100000000: oled_data = 16'b1111011111011110;
				14'b10010110000000: oled_data = 16'b1110011101111110;
				14'b10011000000000: oled_data = 16'b1101111101011101;
				14'b10011010000000: oled_data = 16'b1100011010111100;
				14'b10011100000000: oled_data = 16'b1100011010111100;
				14'b10011110000000: oled_data = 16'b1101011100011101;
				14'b10100000000000: oled_data = 16'b1101011100011101;
				14'b10100010000000: oled_data = 16'b1101111100111101;
				14'b10100100000000: oled_data = 16'b1111011110111110;
				14'b10100110000000: oled_data = 16'b1111111111111111;
				14'b10101000000000: oled_data = 16'b1111111111111111;
				14'b10101010000000: oled_data = 16'b1111111111111111;
				14'b10101100000000: oled_data = 16'b1111111111111111;
				14'b10101110000000: oled_data = 16'b1111111111111111;
				14'b10110000000000: oled_data = 16'b1111111111111111;
				14'b10110010000000: oled_data = 16'b1111111111111111;
				14'b10110100000000: oled_data = 16'b1111111111111111;
				14'b10110110000000: oled_data = 16'b1111111111111111;
				14'b10111000000000: oled_data = 16'b1111111111111111;
				14'b10111010000000: oled_data = 16'b1111111111111111;
				14'b10111100000000: oled_data = 16'b1111111111111111;
				14'b10111110000000: oled_data = 16'b1111111111111111;
				14'b00000000000001: oled_data = 16'b1111111111111111;
				14'b00000010000001: oled_data = 16'b1111111111111111;
				14'b00000100000001: oled_data = 16'b1111111111111111;
				14'b00000110000001: oled_data = 16'b1111111111111111;
				14'b00001000000001: oled_data = 16'b1111111111111111;
				14'b00001010000001: oled_data = 16'b1111111111111111;
				14'b00001100000001: oled_data = 16'b1111111111111111;
				14'b00001110000001: oled_data = 16'b1111111111111111;
				14'b00010000000001: oled_data = 16'b1111111111111111;
				14'b00010010000001: oled_data = 16'b1111111111111111;
				14'b00010100000001: oled_data = 16'b1111111111111111;
				14'b00010110000001: oled_data = 16'b1111111111111111;
				14'b00011000000001: oled_data = 16'b1111111111111111;
				14'b00011010000001: oled_data = 16'b1111111111111111;
				14'b00011100000001: oled_data = 16'b1111111111111111;
				14'b00011110000001: oled_data = 16'b1111111111111111;
				14'b00100000000001: oled_data = 16'b1111111111111111;
				14'b00100010000001: oled_data = 16'b1111111111111111;
				14'b00100100000001: oled_data = 16'b1111111111111111;
				14'b00100110000001: oled_data = 16'b1111111111111111;
				14'b00101000000001: oled_data = 16'b1111111111111111;
				14'b00101010000001: oled_data = 16'b1111111111111111;
				14'b00101100000001: oled_data = 16'b1111111111111111;
				14'b00101110000001: oled_data = 16'b1111111111111111;
				14'b00110000000001: oled_data = 16'b1111111111111111;
				14'b00110010000001: oled_data = 16'b1111111111111111;
				14'b00110100000001: oled_data = 16'b1111111111111111;
				14'b00110110000001: oled_data = 16'b1111111111111111;
				14'b00111000000001: oled_data = 16'b1111111111111111;
				14'b00111010000001: oled_data = 16'b1111111111111111;
				14'b00111100000001: oled_data = 16'b1111111111111111;
				14'b00111110000001: oled_data = 16'b1111111111111111;
				14'b01000000000001: oled_data = 16'b1111111111111111;
				14'b01000010000001: oled_data = 16'b1111111111111111;
				14'b01000100000001: oled_data = 16'b1111111111111111;
				14'b01000110000001: oled_data = 16'b1111111111111111;
				14'b01001000000001: oled_data = 16'b1111111111111111;
				14'b01001010000001: oled_data = 16'b1111111111111111;
				14'b01001100000001: oled_data = 16'b1111111111111111;
				14'b01001110000001: oled_data = 16'b1111111111111111;
				14'b01010000000001: oled_data = 16'b1111111111111111;
				14'b01010010000001: oled_data = 16'b1111111111111111;
				14'b01010100000001: oled_data = 16'b1111111111111111;
				14'b01010110000001: oled_data = 16'b1111111111111111;
				14'b01011000000001: oled_data = 16'b1111111111111111;
				14'b01011010000001: oled_data = 16'b1111111111111111;
				14'b01011100000001: oled_data = 16'b1111111111111111;
				14'b01011110000001: oled_data = 16'b1111111111111111;
				14'b01100000000001: oled_data = 16'b1111111111111111;
				14'b01100010000001: oled_data = 16'b1111111111111111;
				14'b01100100000001: oled_data = 16'b1111111111111111;
				14'b01100110000001: oled_data = 16'b1111111111111111;
				14'b01101000000001: oled_data = 16'b1111111111111111;
				14'b01101010000001: oled_data = 16'b1111111111111111;
				14'b01101100000001: oled_data = 16'b1111111111111111;
				14'b01101110000001: oled_data = 16'b1111111111111111;
				14'b01110000000001: oled_data = 16'b1111111111111111;
				14'b01110010000001: oled_data = 16'b1111111111111111;
				14'b01110100000001: oled_data = 16'b1111111111111111;
				14'b01110110000001: oled_data = 16'b1111111111111111;
				14'b01111000000001: oled_data = 16'b1111111111111111;
				14'b01111010000001: oled_data = 16'b1111111111111111;
				14'b01111100000001: oled_data = 16'b1111111111111111;
				14'b01111110000001: oled_data = 16'b1111111111111111;
				14'b10000000000001: oled_data = 16'b1111111111111111;
				14'b10000010000001: oled_data = 16'b1111111111111111;
				14'b10000100000001: oled_data = 16'b1111111111111111;
				14'b10000110000001: oled_data = 16'b1111111111111111;
				14'b10001000000001: oled_data = 16'b1111111111111111;
				14'b10001010000001: oled_data = 16'b1111111111111111;
				14'b10001100000001: oled_data = 16'b1111111111111111;
				14'b10001110000001: oled_data = 16'b1111111111111111;
				14'b10010000000001: oled_data = 16'b1111111111111111;
				14'b10010010000001: oled_data = 16'b1111111111111111;
				14'b10010100000001: oled_data = 16'b1111011111011110;
				14'b10010110000001: oled_data = 16'b1110011110011110;
				14'b10011000000001: oled_data = 16'b1110011101011101;
				14'b10011010000001: oled_data = 16'b1100111011011100;
				14'b10011100000001: oled_data = 16'b1100011010111100;
				14'b10011110000001: oled_data = 16'b1101011011111101;
				14'b10100000000001: oled_data = 16'b1101011100011101;
				14'b10100010000001: oled_data = 16'b1101111100111101;
				14'b10100100000001: oled_data = 16'b1110111110111110;
				14'b10100110000001: oled_data = 16'b1111111111111111;
				14'b10101000000001: oled_data = 16'b1111111111111111;
				14'b10101010000001: oled_data = 16'b1111111111111111;
				14'b10101100000001: oled_data = 16'b1111111111111111;
				14'b10101110000001: oled_data = 16'b1111111111111111;
				14'b10110000000001: oled_data = 16'b1111111111111111;
				14'b10110010000001: oled_data = 16'b1111111111111111;
				14'b10110100000001: oled_data = 16'b1111111111111111;
				14'b10110110000001: oled_data = 16'b1111111111111111;
				14'b10111000000001: oled_data = 16'b1111111111111111;
				14'b10111010000001: oled_data = 16'b1111111111111111;
				14'b10111100000001: oled_data = 16'b1111111111111111;
				14'b10111110000001: oled_data = 16'b1111111111111111;
				14'b00000000000010: oled_data = 16'b1111111111111111;
				14'b00000010000010: oled_data = 16'b1111111111111111;
				14'b00000100000010: oled_data = 16'b1111111111111111;
				14'b00000110000010: oled_data = 16'b1111111111111111;
				14'b00001000000010: oled_data = 16'b1111111111111111;
				14'b00001010000010: oled_data = 16'b1111111111111111;
				14'b00001100000010: oled_data = 16'b1111111111111111;
				14'b00001110000010: oled_data = 16'b1111111111111111;
				14'b00010000000010: oled_data = 16'b1111111111111111;
				14'b00010010000010: oled_data = 16'b1111111111111111;
				14'b00010100000010: oled_data = 16'b1111111111111111;
				14'b00010110000010: oled_data = 16'b1111111111111111;
				14'b00011000000010: oled_data = 16'b1111111111111111;
				14'b00011010000010: oled_data = 16'b1111111111111111;
				14'b00011100000010: oled_data = 16'b1111111111111111;
				14'b00011110000010: oled_data = 16'b1111111111111111;
				14'b00100000000010: oled_data = 16'b1111111111111111;
				14'b00100010000010: oled_data = 16'b1111111111111111;
				14'b00100100000010: oled_data = 16'b1111111111111111;
				14'b00100110000010: oled_data = 16'b1111111111111111;
				14'b00101000000010: oled_data = 16'b1111111111111111;
				14'b00101010000010: oled_data = 16'b1111111111111111;
				14'b00101100000010: oled_data = 16'b1111111111111111;
				14'b00101110000010: oled_data = 16'b1111111111111111;
				14'b00110000000010: oled_data = 16'b1111111111111111;
				14'b00110010000010: oled_data = 16'b1111111111111111;
				14'b00110100000010: oled_data = 16'b1111111111111111;
				14'b00110110000010: oled_data = 16'b1111111111111111;
				14'b00111000000010: oled_data = 16'b1111111111111111;
				14'b00111010000010: oled_data = 16'b1111111111111111;
				14'b00111100000010: oled_data = 16'b1111111111111111;
				14'b00111110000010: oled_data = 16'b1111111111111111;
				14'b01000000000010: oled_data = 16'b1111111111111111;
				14'b01000010000010: oled_data = 16'b1111111111111111;
				14'b01000100000010: oled_data = 16'b1111111111111111;
				14'b01000110000010: oled_data = 16'b1111111111111111;
				14'b01001000000010: oled_data = 16'b1111111111111111;
				14'b01001010000010: oled_data = 16'b1111111111111111;
				14'b01001100000010: oled_data = 16'b1111111111111111;
				14'b01001110000010: oled_data = 16'b1111111111111111;
				14'b01010000000010: oled_data = 16'b1111111111111111;
				14'b01010010000010: oled_data = 16'b1111111111111111;
				14'b01010100000010: oled_data = 16'b1111111111111111;
				14'b01010110000010: oled_data = 16'b1111111111111111;
				14'b01011000000010: oled_data = 16'b1111111111111111;
				14'b01011010000010: oled_data = 16'b1111111111111111;
				14'b01011100000010: oled_data = 16'b1111111111111111;
				14'b01011110000010: oled_data = 16'b1111111111111111;
				14'b01100000000010: oled_data = 16'b1111111111111111;
				14'b01100010000010: oled_data = 16'b1111111111111111;
				14'b01100100000010: oled_data = 16'b1111111111111111;
				14'b01100110000010: oled_data = 16'b1111111111111111;
				14'b01101000000010: oled_data = 16'b1111111111111111;
				14'b01101010000010: oled_data = 16'b1111111111111111;
				14'b01101100000010: oled_data = 16'b1111111111111111;
				14'b01101110000010: oled_data = 16'b1111111111111111;
				14'b01110000000010: oled_data = 16'b1111111111111111;
				14'b01110010000010: oled_data = 16'b1111111111111111;
				14'b01110100000010: oled_data = 16'b1111111111111111;
				14'b01110110000010: oled_data = 16'b1111111111111111;
				14'b01111000000010: oled_data = 16'b1111111111111111;
				14'b01111010000010: oled_data = 16'b1111111111111111;
				14'b01111100000010: oled_data = 16'b1111111111111111;
				14'b01111110000010: oled_data = 16'b1111111111111111;
				14'b10000000000010: oled_data = 16'b1111111111111111;
				14'b10000010000010: oled_data = 16'b1111111111111111;
				14'b10000100000010: oled_data = 16'b1111111111111111;
				14'b10000110000010: oled_data = 16'b1111111111111111;
				14'b10001000000010: oled_data = 16'b1111111111111111;
				14'b10001010000010: oled_data = 16'b1111111111111111;
				14'b10001100000010: oled_data = 16'b1111111111111111;
				14'b10001110000010: oled_data = 16'b1111111111111111;
				14'b10010000000010: oled_data = 16'b1111111111111111;
				14'b10010010000010: oled_data = 16'b1111111111111111;
				14'b10010100000010: oled_data = 16'b1111011111011110;
				14'b10010110000010: oled_data = 16'b1110111110011110;
				14'b10011000000010: oled_data = 16'b1110011101111101;
				14'b10011010000010: oled_data = 16'b1100111011111100;
				14'b10011100000010: oled_data = 16'b1100011011011100;
				14'b10011110000010: oled_data = 16'b1101011011111100;
				14'b10100000000010: oled_data = 16'b1101011100011101;
				14'b10100010000010: oled_data = 16'b1101011100011101;
				14'b10100100000010: oled_data = 16'b1110111110011110;
				14'b10100110000010: oled_data = 16'b1111111111111111;
				14'b10101000000010: oled_data = 16'b1111111111111111;
				14'b10101010000010: oled_data = 16'b1111111111111111;
				14'b10101100000010: oled_data = 16'b1111111111111111;
				14'b10101110000010: oled_data = 16'b1111111111111111;
				14'b10110000000010: oled_data = 16'b1111111111111111;
				14'b10110010000010: oled_data = 16'b1111111111111111;
				14'b10110100000010: oled_data = 16'b1111111111111111;
				14'b10110110000010: oled_data = 16'b1111111111111111;
				14'b10111000000010: oled_data = 16'b1111111111111111;
				14'b10111010000010: oled_data = 16'b1111111111111111;
				14'b10111100000010: oled_data = 16'b1111111111111111;
				14'b10111110000010: oled_data = 16'b1111111111111111;
				14'b00000000000011: oled_data = 16'b1111111111111111;
				14'b00000010000011: oled_data = 16'b1111111111111111;
				14'b00000100000011: oled_data = 16'b1111111111111111;
				14'b00000110000011: oled_data = 16'b1111111111111111;
				14'b00001000000011: oled_data = 16'b1111111111111111;
				14'b00001010000011: oled_data = 16'b1111111111111111;
				14'b00001100000011: oled_data = 16'b1111111111111111;
				14'b00001110000011: oled_data = 16'b1111111111111111;
				14'b00010000000011: oled_data = 16'b1111111111111111;
				14'b00010010000011: oled_data = 16'b1111111111111111;
				14'b00010100000011: oled_data = 16'b1111111111111111;
				14'b00010110000011: oled_data = 16'b1111111111111111;
				14'b00011000000011: oled_data = 16'b1111111111111111;
				14'b00011010000011: oled_data = 16'b1111111111111111;
				14'b00011100000011: oled_data = 16'b1111111111111111;
				14'b00011110000011: oled_data = 16'b1111111111111111;
				14'b00100000000011: oled_data = 16'b1111111111111111;
				14'b00100010000011: oled_data = 16'b1111111111111111;
				14'b00100100000011: oled_data = 16'b1111111111111111;
				14'b00100110000011: oled_data = 16'b1111111111111111;
				14'b00101000000011: oled_data = 16'b1111111111111111;
				14'b00101010000011: oled_data = 16'b1111111111111111;
				14'b00101100000011: oled_data = 16'b1111111111111111;
				14'b00101110000011: oled_data = 16'b1111111111111111;
				14'b00110000000011: oled_data = 16'b1111111111111111;
				14'b00110010000011: oled_data = 16'b1111111111111111;
				14'b00110100000011: oled_data = 16'b1111111111111111;
				14'b00110110000011: oled_data = 16'b1111111111111111;
				14'b00111000000011: oled_data = 16'b1111111111111111;
				14'b00111010000011: oled_data = 16'b1111111111111111;
				14'b00111100000011: oled_data = 16'b1111111111111111;
				14'b00111110000011: oled_data = 16'b1111111111111111;
				14'b01000000000011: oled_data = 16'b1111111111111111;
				14'b01000010000011: oled_data = 16'b1111111111111111;
				14'b01000100000011: oled_data = 16'b1111111111111111;
				14'b01000110000011: oled_data = 16'b1111111111111111;
				14'b01001000000011: oled_data = 16'b1111111111111111;
				14'b01001010000011: oled_data = 16'b1111111111111111;
				14'b01001100000011: oled_data = 16'b1111111111111111;
				14'b01001110000011: oled_data = 16'b1111111111111111;
				14'b01010000000011: oled_data = 16'b1111111111111111;
				14'b01010010000011: oled_data = 16'b1111111111111111;
				14'b01010100000011: oled_data = 16'b1111111111111111;
				14'b01010110000011: oled_data = 16'b1111111111111111;
				14'b01011000000011: oled_data = 16'b1111111111111111;
				14'b01011010000011: oled_data = 16'b1111111111111111;
				14'b01011100000011: oled_data = 16'b1111111111111111;
				14'b01011110000011: oled_data = 16'b1111111111111111;
				14'b01100000000011: oled_data = 16'b1111111111111111;
				14'b01100010000011: oled_data = 16'b1111111111111111;
				14'b01100100000011: oled_data = 16'b1111111111111111;
				14'b01100110000011: oled_data = 16'b1111111111111111;
				14'b01101000000011: oled_data = 16'b1111111111111111;
				14'b01101010000011: oled_data = 16'b1111111111111111;
				14'b01101100000011: oled_data = 16'b1111111111111111;
				14'b01101110000011: oled_data = 16'b1111111111111111;
				14'b01110000000011: oled_data = 16'b1111111111111111;
				14'b01110010000011: oled_data = 16'b1111111111111111;
				14'b01110100000011: oled_data = 16'b1111111111111111;
				14'b01110110000011: oled_data = 16'b1111111111111111;
				14'b01111000000011: oled_data = 16'b1111111111111111;
				14'b01111010000011: oled_data = 16'b1111111111111111;
				14'b01111100000011: oled_data = 16'b1111111111111111;
				14'b01111110000011: oled_data = 16'b1111111111111111;
				14'b10000000000011: oled_data = 16'b1111111111111111;
				14'b10000010000011: oled_data = 16'b1111111111111111;
				14'b10000100000011: oled_data = 16'b1111111111111111;
				14'b10000110000011: oled_data = 16'b1111111111111111;
				14'b10001000000011: oled_data = 16'b1111111111111111;
				14'b10001010000011: oled_data = 16'b1111111111111111;
				14'b10001100000011: oled_data = 16'b1111111111111111;
				14'b10001110000011: oled_data = 16'b1111111111111111;
				14'b10010000000011: oled_data = 16'b1111111111111111;
				14'b10010010000011: oled_data = 16'b1111111111111111;
				14'b10010100000011: oled_data = 16'b1111111111111111;
				14'b10010110000011: oled_data = 16'b1110111110011110;
				14'b10011000000011: oled_data = 16'b1110011101111101;
				14'b10011010000011: oled_data = 16'b1101011100011100;
				14'b10011100000011: oled_data = 16'b1100011011011100;
				14'b10011110000011: oled_data = 16'b1100111011111100;
				14'b10100000000011: oled_data = 16'b1101011100011101;
				14'b10100010000011: oled_data = 16'b1101011100011101;
				14'b10100100000011: oled_data = 16'b1110011101111101;
				14'b10100110000011: oled_data = 16'b1111011111011110;
				14'b10101000000011: oled_data = 16'b1111111111111111;
				14'b10101010000011: oled_data = 16'b1111111111111111;
				14'b10101100000011: oled_data = 16'b1111111111111111;
				14'b10101110000011: oled_data = 16'b1111111111111111;
				14'b10110000000011: oled_data = 16'b1111111111111111;
				14'b10110010000011: oled_data = 16'b1111111111111111;
				14'b10110100000011: oled_data = 16'b1111111111111111;
				14'b10110110000011: oled_data = 16'b1111111111111111;
				14'b10111000000011: oled_data = 16'b1111111111111111;
				14'b10111010000011: oled_data = 16'b1111111111111111;
				14'b10111100000011: oled_data = 16'b1111111111111111;
				14'b10111110000011: oled_data = 16'b1111111111111111;
				14'b00000000000100: oled_data = 16'b1111111111111111;
				14'b00000010000100: oled_data = 16'b1111111111111111;
				14'b00000100000100: oled_data = 16'b1111111111111111;
				14'b00000110000100: oled_data = 16'b1111111111111111;
				14'b00001000000100: oled_data = 16'b1111111111111111;
				14'b00001010000100: oled_data = 16'b1111111111111111;
				14'b00001100000100: oled_data = 16'b1111111111111111;
				14'b00001110000100: oled_data = 16'b1111111111111111;
				14'b00010000000100: oled_data = 16'b1111111111111111;
				14'b00010010000100: oled_data = 16'b1111111111111111;
				14'b00010100000100: oled_data = 16'b1111111111111111;
				14'b00010110000100: oled_data = 16'b1111111111111111;
				14'b00011000000100: oled_data = 16'b1111111111111111;
				14'b00011010000100: oled_data = 16'b1111111111111111;
				14'b00011100000100: oled_data = 16'b1111111111111111;
				14'b00011110000100: oled_data = 16'b1111111111111111;
				14'b00100000000100: oled_data = 16'b1111111111111111;
				14'b00100010000100: oled_data = 16'b1111111111111111;
				14'b00100100000100: oled_data = 16'b1111111111111111;
				14'b00100110000100: oled_data = 16'b1111111111111111;
				14'b00101000000100: oled_data = 16'b1111111111111111;
				14'b00101010000100: oled_data = 16'b1111111111111111;
				14'b00101100000100: oled_data = 16'b1111111111111111;
				14'b00101110000100: oled_data = 16'b1111111111111111;
				14'b00110000000100: oled_data = 16'b1111111111111111;
				14'b00110010000100: oled_data = 16'b1111111111111111;
				14'b00110100000100: oled_data = 16'b1111111111111111;
				14'b00110110000100: oled_data = 16'b1111111111111111;
				14'b00111000000100: oled_data = 16'b1111111111111111;
				14'b00111010000100: oled_data = 16'b1111111111111111;
				14'b00111100000100: oled_data = 16'b1111111111111111;
				14'b00111110000100: oled_data = 16'b1111111111111111;
				14'b01000000000100: oled_data = 16'b1111111111111111;
				14'b01000010000100: oled_data = 16'b1111111111111111;
				14'b01000100000100: oled_data = 16'b1111111111111111;
				14'b01000110000100: oled_data = 16'b1111111111111111;
				14'b01001000000100: oled_data = 16'b1111111111111111;
				14'b01001010000100: oled_data = 16'b1111111111111111;
				14'b01001100000100: oled_data = 16'b1111111111111111;
				14'b01001110000100: oled_data = 16'b1111111111111111;
				14'b01010000000100: oled_data = 16'b1111111111111111;
				14'b01010010000100: oled_data = 16'b1111111111111111;
				14'b01010100000100: oled_data = 16'b1111111111111111;
				14'b01010110000100: oled_data = 16'b1111111111111111;
				14'b01011000000100: oled_data = 16'b1111111111111111;
				14'b01011010000100: oled_data = 16'b1111111111111111;
				14'b01011100000100: oled_data = 16'b1111111111111111;
				14'b01011110000100: oled_data = 16'b1111111111111111;
				14'b01100000000100: oled_data = 16'b1111111111111111;
				14'b01100010000100: oled_data = 16'b1111111111111111;
				14'b01100100000100: oled_data = 16'b1111111111111111;
				14'b01100110000100: oled_data = 16'b1111111111111111;
				14'b01101000000100: oled_data = 16'b1111111111111111;
				14'b01101010000100: oled_data = 16'b1111111111111111;
				14'b01101100000100: oled_data = 16'b1111111111111111;
				14'b01101110000100: oled_data = 16'b1111111111111111;
				14'b01110000000100: oled_data = 16'b1111111111111111;
				14'b01110010000100: oled_data = 16'b1111111111111111;
				14'b01110100000100: oled_data = 16'b1111111111111111;
				14'b01110110000100: oled_data = 16'b1111111111111111;
				14'b01111000000100: oled_data = 16'b1111111111111111;
				14'b01111010000100: oled_data = 16'b1111111111111111;
				14'b01111100000100: oled_data = 16'b1111111111111111;
				14'b01111110000100: oled_data = 16'b1111111111111111;
				14'b10000000000100: oled_data = 16'b1111111111111111;
				14'b10000010000100: oled_data = 16'b1111111111111111;
				14'b10000100000100: oled_data = 16'b1111111111111111;
				14'b10000110000100: oled_data = 16'b1111111111111111;
				14'b10001000000100: oled_data = 16'b1111111111111111;
				14'b10001010000100: oled_data = 16'b1111111111111111;
				14'b10001100000100: oled_data = 16'b1111111111111111;
				14'b10001110000100: oled_data = 16'b1111111111111111;
				14'b10010000000100: oled_data = 16'b1111111111111111;
				14'b10010010000100: oled_data = 16'b1111111111111111;
				14'b10010100000100: oled_data = 16'b1111111111111111;
				14'b10010110000100: oled_data = 16'b1110111110111110;
				14'b10011000000100: oled_data = 16'b1110011101111101;
				14'b10011010000100: oled_data = 16'b1101011100111101;
				14'b10011100000100: oled_data = 16'b1100011011011011;
				14'b10011110000100: oled_data = 16'b1100111011011100;
				14'b10100000000100: oled_data = 16'b1101011100011100;
				14'b10100010000100: oled_data = 16'b1101011100011100;
				14'b10100100000100: oled_data = 16'b1101111101011101;
				14'b10100110000100: oled_data = 16'b1111011111011110;
				14'b10101000000100: oled_data = 16'b1111111111111111;
				14'b10101010000100: oled_data = 16'b1111111111111111;
				14'b10101100000100: oled_data = 16'b1111111111111111;
				14'b10101110000100: oled_data = 16'b1111111111111111;
				14'b10110000000100: oled_data = 16'b1111111111111111;
				14'b10110010000100: oled_data = 16'b1111111111111111;
				14'b10110100000100: oled_data = 16'b1111111111111111;
				14'b10110110000100: oled_data = 16'b1111111111111111;
				14'b10111000000100: oled_data = 16'b1111111111111111;
				14'b10111010000100: oled_data = 16'b1111111111111111;
				14'b10111100000100: oled_data = 16'b1111111111111111;
				14'b10111110000100: oled_data = 16'b1111111111111111;
				14'b00000000000101: oled_data = 16'b1111111111111111;
				14'b00000010000101: oled_data = 16'b1111111111111111;
				14'b00000100000101: oled_data = 16'b1111111111111111;
				14'b00000110000101: oled_data = 16'b1111111111111111;
				14'b00001000000101: oled_data = 16'b1111111111111111;
				14'b00001010000101: oled_data = 16'b1111111111111111;
				14'b00001100000101: oled_data = 16'b1111111111111111;
				14'b00001110000101: oled_data = 16'b1111111111111111;
				14'b00010000000101: oled_data = 16'b1111111111111111;
				14'b00010010000101: oled_data = 16'b1111111111111111;
				14'b00010100000101: oled_data = 16'b1111111111111111;
				14'b00010110000101: oled_data = 16'b1111111111111111;
				14'b00011000000101: oled_data = 16'b1111111111111111;
				14'b00011010000101: oled_data = 16'b1111111111111111;
				14'b00011100000101: oled_data = 16'b1111111111111111;
				14'b00011110000101: oled_data = 16'b1111111111111111;
				14'b00100000000101: oled_data = 16'b1111111111111111;
				14'b00100010000101: oled_data = 16'b1111111111111111;
				14'b00100100000101: oled_data = 16'b1111111111111111;
				14'b00100110000101: oled_data = 16'b1111111111111111;
				14'b00101000000101: oled_data = 16'b1111111111111111;
				14'b00101010000101: oled_data = 16'b1111111111111111;
				14'b00101100000101: oled_data = 16'b1111111111111111;
				14'b00101110000101: oled_data = 16'b1111111111111111;
				14'b00110000000101: oled_data = 16'b1111111111111111;
				14'b00110010000101: oled_data = 16'b1111111111111111;
				14'b00110100000101: oled_data = 16'b1111111111111111;
				14'b00110110000101: oled_data = 16'b1111111111111111;
				14'b00111000000101: oled_data = 16'b1111111111111111;
				14'b00111010000101: oled_data = 16'b1111111111111111;
				14'b00111100000101: oled_data = 16'b1111111111111111;
				14'b00111110000101: oled_data = 16'b1111111111111111;
				14'b01000000000101: oled_data = 16'b1111111111111111;
				14'b01000010000101: oled_data = 16'b1111111111111111;
				14'b01000100000101: oled_data = 16'b1111111111111111;
				14'b01000110000101: oled_data = 16'b1111111111111111;
				14'b01001000000101: oled_data = 16'b1111111111111111;
				14'b01001010000101: oled_data = 16'b1111111111111111;
				14'b01001100000101: oled_data = 16'b1111111111111111;
				14'b01001110000101: oled_data = 16'b1111111111111111;
				14'b01010000000101: oled_data = 16'b1111111111111111;
				14'b01010010000101: oled_data = 16'b1111111111111111;
				14'b01010100000101: oled_data = 16'b1111111111111111;
				14'b01010110000101: oled_data = 16'b1111111111111111;
				14'b01011000000101: oled_data = 16'b1111111111111111;
				14'b01011010000101: oled_data = 16'b1111111111111111;
				14'b01011100000101: oled_data = 16'b1111111111111111;
				14'b01011110000101: oled_data = 16'b1111111111111111;
				14'b01100000000101: oled_data = 16'b1111111111111111;
				14'b01100010000101: oled_data = 16'b1111111111111111;
				14'b01100100000101: oled_data = 16'b1111111111111111;
				14'b01100110000101: oled_data = 16'b1111111111111111;
				14'b01101000000101: oled_data = 16'b1111111111111111;
				14'b01101010000101: oled_data = 16'b1111111111111111;
				14'b01101100000101: oled_data = 16'b1111111111111111;
				14'b01101110000101: oled_data = 16'b1111111111111111;
				14'b01110000000101: oled_data = 16'b1111111111111111;
				14'b01110010000101: oled_data = 16'b1111111111111111;
				14'b01110100000101: oled_data = 16'b1111111111111111;
				14'b01110110000101: oled_data = 16'b1111111111111111;
				14'b01111000000101: oled_data = 16'b1111111111111111;
				14'b01111010000101: oled_data = 16'b1111111111111111;
				14'b01111100000101: oled_data = 16'b1111111111111111;
				14'b01111110000101: oled_data = 16'b1111111111111111;
				14'b10000000000101: oled_data = 16'b1111111111111111;
				14'b10000010000101: oled_data = 16'b1111111111111111;
				14'b10000100000101: oled_data = 16'b1111111111111111;
				14'b10000110000101: oled_data = 16'b1111111111111111;
				14'b10001000000101: oled_data = 16'b1111111111111111;
				14'b10001010000101: oled_data = 16'b1111111111111111;
				14'b10001100000101: oled_data = 16'b1111111111111111;
				14'b10001110000101: oled_data = 16'b1111111111111111;
				14'b10010000000101: oled_data = 16'b1111111111111111;
				14'b10010010000101: oled_data = 16'b1111111111111111;
				14'b10010100000101: oled_data = 16'b1111111111111111;
				14'b10010110000101: oled_data = 16'b1111011111011110;
				14'b10011000000101: oled_data = 16'b1110011101111101;
				14'b10011010000101: oled_data = 16'b1101111101011101;
				14'b10011100000101: oled_data = 16'b1100011011011011;
				14'b10011110000101: oled_data = 16'b1100111011011011;
				14'b10100000000101: oled_data = 16'b1101011100011100;
				14'b10100010000101: oled_data = 16'b1101011100011100;
				14'b10100100000101: oled_data = 16'b1101111100111101;
				14'b10100110000101: oled_data = 16'b1110111110111110;
				14'b10101000000101: oled_data = 16'b1111111111111111;
				14'b10101010000101: oled_data = 16'b1111111111111111;
				14'b10101100000101: oled_data = 16'b1111111111111111;
				14'b10101110000101: oled_data = 16'b1111111111111111;
				14'b10110000000101: oled_data = 16'b1111111111111111;
				14'b10110010000101: oled_data = 16'b1111111111111111;
				14'b10110100000101: oled_data = 16'b1111111111111111;
				14'b10110110000101: oled_data = 16'b1111111111111111;
				14'b10111000000101: oled_data = 16'b1111111111111111;
				14'b10111010000101: oled_data = 16'b1111111111111111;
				14'b10111100000101: oled_data = 16'b1111111111111111;
				14'b10111110000101: oled_data = 16'b1111111111111111;
				14'b00000000000110: oled_data = 16'b1111111111111111;
				14'b00000010000110: oled_data = 16'b1111111111111111;
				14'b00000100000110: oled_data = 16'b1111111111111111;
				14'b00000110000110: oled_data = 16'b1111111111111111;
				14'b00001000000110: oled_data = 16'b1111111111111111;
				14'b00001010000110: oled_data = 16'b1111111111111111;
				14'b00001100000110: oled_data = 16'b1111111111111111;
				14'b00001110000110: oled_data = 16'b1111111111111111;
				14'b00010000000110: oled_data = 16'b1111111111111111;
				14'b00010010000110: oled_data = 16'b1111111111111111;
				14'b00010100000110: oled_data = 16'b1111111111111111;
				14'b00010110000110: oled_data = 16'b1111111111111111;
				14'b00011000000110: oled_data = 16'b1111111111111111;
				14'b00011010000110: oled_data = 16'b1111111111111111;
				14'b00011100000110: oled_data = 16'b1111111111111111;
				14'b00011110000110: oled_data = 16'b1111111111111111;
				14'b00100000000110: oled_data = 16'b1111111111111111;
				14'b00100010000110: oled_data = 16'b1111111111111111;
				14'b00100100000110: oled_data = 16'b1111111111111111;
				14'b00100110000110: oled_data = 16'b1111111111111111;
				14'b00101000000110: oled_data = 16'b1111111111111111;
				14'b00101010000110: oled_data = 16'b1111111111111111;
				14'b00101100000110: oled_data = 16'b1111111111111111;
				14'b00101110000110: oled_data = 16'b1111111111111111;
				14'b00110000000110: oled_data = 16'b1111111111111111;
				14'b00110010000110: oled_data = 16'b1111111111111111;
				14'b00110100000110: oled_data = 16'b1111111111111111;
				14'b00110110000110: oled_data = 16'b1111111111111111;
				14'b00111000000110: oled_data = 16'b1111111111111111;
				14'b00111010000110: oled_data = 16'b1111111111111111;
				14'b00111100000110: oled_data = 16'b1111111111111111;
				14'b00111110000110: oled_data = 16'b1111111111111111;
				14'b01000000000110: oled_data = 16'b1111111111111111;
				14'b01000010000110: oled_data = 16'b1111111111111111;
				14'b01000100000110: oled_data = 16'b1111111111111111;
				14'b01000110000110: oled_data = 16'b1111111111111111;
				14'b01001000000110: oled_data = 16'b1111111111111111;
				14'b01001010000110: oled_data = 16'b1111111111111111;
				14'b01001100000110: oled_data = 16'b1111111111111111;
				14'b01001110000110: oled_data = 16'b1111111111111111;
				14'b01010000000110: oled_data = 16'b1111111111111111;
				14'b01010010000110: oled_data = 16'b1111111111111111;
				14'b01010100000110: oled_data = 16'b1111111111111111;
				14'b01010110000110: oled_data = 16'b1111111111111111;
				14'b01011000000110: oled_data = 16'b1111111111111111;
				14'b01011010000110: oled_data = 16'b1111111111111111;
				14'b01011100000110: oled_data = 16'b1111111111111111;
				14'b01011110000110: oled_data = 16'b1111111111111111;
				14'b01100000000110: oled_data = 16'b1111111111111111;
				14'b01100010000110: oled_data = 16'b1111111111111111;
				14'b01100100000110: oled_data = 16'b1111111111111111;
				14'b01100110000110: oled_data = 16'b1111111111111111;
				14'b01101000000110: oled_data = 16'b1111111111111111;
				14'b01101010000110: oled_data = 16'b1111111111111111;
				14'b01101100000110: oled_data = 16'b1111111111111111;
				14'b01101110000110: oled_data = 16'b1111111111111111;
				14'b01110000000110: oled_data = 16'b1111111111111111;
				14'b01110010000110: oled_data = 16'b1111111111111111;
				14'b01110100000110: oled_data = 16'b1111111111111111;
				14'b01110110000110: oled_data = 16'b1111111111111111;
				14'b01111000000110: oled_data = 16'b1111111111111111;
				14'b01111010000110: oled_data = 16'b1111111111111111;
				14'b01111100000110: oled_data = 16'b1111111111111111;
				14'b01111110000110: oled_data = 16'b1111111111111111;
				14'b10000000000110: oled_data = 16'b1111111111111111;
				14'b10000010000110: oled_data = 16'b1111111111111111;
				14'b10000100000110: oled_data = 16'b1111111111111111;
				14'b10000110000110: oled_data = 16'b1111111111111111;
				14'b10001000000110: oled_data = 16'b1111111111111111;
				14'b10001010000110: oled_data = 16'b1111111111111111;
				14'b10001100000110: oled_data = 16'b1111111111111111;
				14'b10001110000110: oled_data = 16'b1111111111111111;
				14'b10010000000110: oled_data = 16'b1111111111111111;
				14'b10010010000110: oled_data = 16'b1111111111111111;
				14'b10010100000110: oled_data = 16'b1111111111111111;
				14'b10010110000110: oled_data = 16'b1111011111011110;
				14'b10011000000110: oled_data = 16'b1110011110011101;
				14'b10011010000110: oled_data = 16'b1110011101111101;
				14'b10011100000110: oled_data = 16'b1100111011111011;
				14'b10011110000110: oled_data = 16'b1100011011011011;
				14'b10100000000110: oled_data = 16'b1101011011111100;
				14'b10100010000110: oled_data = 16'b1101011100011100;
				14'b10100100000110: oled_data = 16'b1101011100011100;
				14'b10100110000110: oled_data = 16'b1110011101111101;
				14'b10101000000110: oled_data = 16'b1111011111011110;
				14'b10101010000110: oled_data = 16'b1111111111111111;
				14'b10101100000110: oled_data = 16'b1111111111111111;
				14'b10101110000110: oled_data = 16'b1111111111111111;
				14'b10110000000110: oled_data = 16'b1111111111111111;
				14'b10110010000110: oled_data = 16'b1111111111111111;
				14'b10110100000110: oled_data = 16'b1111111111111111;
				14'b10110110000110: oled_data = 16'b1111111111111111;
				14'b10111000000110: oled_data = 16'b1111111111111111;
				14'b10111010000110: oled_data = 16'b1111111111111111;
				14'b10111100000110: oled_data = 16'b1111111111111111;
				14'b10111110000110: oled_data = 16'b1111111111111111;
				14'b00000000000111: oled_data = 16'b1111111111111111;
				14'b00000010000111: oled_data = 16'b1111111111111111;
				14'b00000100000111: oled_data = 16'b1111111111111111;
				14'b00000110000111: oled_data = 16'b1111111111111111;
				14'b00001000000111: oled_data = 16'b1111111111111111;
				14'b00001010000111: oled_data = 16'b1111111111111111;
				14'b00001100000111: oled_data = 16'b1111111111111111;
				14'b00001110000111: oled_data = 16'b1111111111111111;
				14'b00010000000111: oled_data = 16'b1111111111111111;
				14'b00010010000111: oled_data = 16'b1111111111111111;
				14'b00010100000111: oled_data = 16'b1111111111111111;
				14'b00010110000111: oled_data = 16'b1111111111111111;
				14'b00011000000111: oled_data = 16'b1111111111111111;
				14'b00011010000111: oled_data = 16'b1111111111111111;
				14'b00011100000111: oled_data = 16'b1111111111111111;
				14'b00011110000111: oled_data = 16'b1111111111111111;
				14'b00100000000111: oled_data = 16'b1111111111111111;
				14'b00100010000111: oled_data = 16'b1111111111111111;
				14'b00100100000111: oled_data = 16'b1111111111111111;
				14'b00100110000111: oled_data = 16'b1111111111111111;
				14'b00101000000111: oled_data = 16'b1111111111111111;
				14'b00101010000111: oled_data = 16'b1111111111111111;
				14'b00101100000111: oled_data = 16'b1111111111111111;
				14'b00101110000111: oled_data = 16'b1111111111111111;
				14'b00110000000111: oled_data = 16'b1111111111111111;
				14'b00110010000111: oled_data = 16'b1111111111111111;
				14'b00110100000111: oled_data = 16'b1111111111111111;
				14'b00110110000111: oled_data = 16'b1111111111111111;
				14'b00111000000111: oled_data = 16'b1111111111111111;
				14'b00111010000111: oled_data = 16'b1111111111111111;
				14'b00111100000111: oled_data = 16'b1111111111111111;
				14'b00111110000111: oled_data = 16'b1111111111111111;
				14'b01000000000111: oled_data = 16'b1111111111111111;
				14'b01000010000111: oled_data = 16'b1111111111111111;
				14'b01000100000111: oled_data = 16'b1111111111111111;
				14'b01000110000111: oled_data = 16'b1111111111111111;
				14'b01001000000111: oled_data = 16'b1111111111111111;
				14'b01001010000111: oled_data = 16'b1111111111111111;
				14'b01001100000111: oled_data = 16'b1111111111111111;
				14'b01001110000111: oled_data = 16'b1111111111111111;
				14'b01010000000111: oled_data = 16'b1111111111111111;
				14'b01010010000111: oled_data = 16'b1111111111111111;
				14'b01010100000111: oled_data = 16'b1111111111111111;
				14'b01010110000111: oled_data = 16'b1111111111111111;
				14'b01011000000111: oled_data = 16'b1111111111111111;
				14'b01011010000111: oled_data = 16'b1111111111111111;
				14'b01011100000111: oled_data = 16'b1111111111111111;
				14'b01011110000111: oled_data = 16'b1111111111111111;
				14'b01100000000111: oled_data = 16'b1111111111111111;
				14'b01100010000111: oled_data = 16'b1111111111111111;
				14'b01100100000111: oled_data = 16'b1111111111111111;
				14'b01100110000111: oled_data = 16'b1111111111111111;
				14'b01101000000111: oled_data = 16'b1111111111111111;
				14'b01101010000111: oled_data = 16'b1111111111111111;
				14'b01101100000111: oled_data = 16'b1111111111111111;
				14'b01101110000111: oled_data = 16'b1111111111111111;
				14'b01110000000111: oled_data = 16'b1111111111111111;
				14'b01110010000111: oled_data = 16'b1111111111111111;
				14'b01110100000111: oled_data = 16'b1111111111111111;
				14'b01110110000111: oled_data = 16'b1111111111111111;
				14'b01111000000111: oled_data = 16'b1111111111111111;
				14'b01111010000111: oled_data = 16'b1111111111111111;
				14'b01111100000111: oled_data = 16'b1111111111111111;
				14'b01111110000111: oled_data = 16'b1111111111111111;
				14'b10000000000111: oled_data = 16'b1111111111111111;
				14'b10000010000111: oled_data = 16'b1111111111111111;
				14'b10000100000111: oled_data = 16'b1111111111111111;
				14'b10000110000111: oled_data = 16'b1111111111111111;
				14'b10001000000111: oled_data = 16'b1111111111111111;
				14'b10001010000111: oled_data = 16'b1111111111111111;
				14'b10001100000111: oled_data = 16'b1111111111111111;
				14'b10001110000111: oled_data = 16'b1111111111111111;
				14'b10010000000111: oled_data = 16'b1111111111111111;
				14'b10010010000111: oled_data = 16'b1111111111111111;
				14'b10010100000111: oled_data = 16'b1111111111111111;
				14'b10010110000111: oled_data = 16'b1111111111111111;
				14'b10011000000111: oled_data = 16'b1110111110011110;
				14'b10011010000111: oled_data = 16'b1110011110011101;
				14'b10011100000111: oled_data = 16'b1101011100011100;
				14'b10011110000111: oled_data = 16'b1100011011011011;
				14'b10100000000111: oled_data = 16'b1100111011111011;
				14'b10100010000111: oled_data = 16'b1101011100111100;
				14'b10100100000111: oled_data = 16'b1101011100011100;
				14'b10100110000111: oled_data = 16'b1101111101011101;
				14'b10101000000111: oled_data = 16'b1111011110111110;
				14'b10101010000111: oled_data = 16'b1111111111111111;
				14'b10101100000111: oled_data = 16'b1111111111111111;
				14'b10101110000111: oled_data = 16'b1111111111111111;
				14'b10110000000111: oled_data = 16'b1111111111111111;
				14'b10110010000111: oled_data = 16'b1111111111111111;
				14'b10110100000111: oled_data = 16'b1111111111111111;
				14'b10110110000111: oled_data = 16'b1111111111111111;
				14'b10111000000111: oled_data = 16'b1111111111111111;
				14'b10111010000111: oled_data = 16'b1111111111111111;
				14'b10111100000111: oled_data = 16'b1111111111111111;
				14'b10111110000111: oled_data = 16'b1111111111111111;
				14'b00000000001000: oled_data = 16'b1111111111111111;
				14'b00000010001000: oled_data = 16'b1111111111111111;
				14'b00000100001000: oled_data = 16'b1111111111111111;
				14'b00000110001000: oled_data = 16'b1111111111111111;
				14'b00001000001000: oled_data = 16'b1111111111111111;
				14'b00001010001000: oled_data = 16'b1111111111111111;
				14'b00001100001000: oled_data = 16'b1111111111111111;
				14'b00001110001000: oled_data = 16'b1111111111111111;
				14'b00010000001000: oled_data = 16'b1111111111111111;
				14'b00010010001000: oled_data = 16'b1111111111111111;
				14'b00010100001000: oled_data = 16'b1111111111111111;
				14'b00010110001000: oled_data = 16'b1111111111111111;
				14'b00011000001000: oled_data = 16'b1111111111111111;
				14'b00011010001000: oled_data = 16'b1111111111111111;
				14'b00011100001000: oled_data = 16'b1111111111111111;
				14'b00011110001000: oled_data = 16'b1111111111111111;
				14'b00100000001000: oled_data = 16'b1111111111111111;
				14'b00100010001000: oled_data = 16'b1111111111111111;
				14'b00100100001000: oled_data = 16'b1111111111111111;
				14'b00100110001000: oled_data = 16'b1111111111111111;
				14'b00101000001000: oled_data = 16'b1111111111111111;
				14'b00101010001000: oled_data = 16'b1111111111111111;
				14'b00101100001000: oled_data = 16'b1111111111111111;
				14'b00101110001000: oled_data = 16'b1111111111111111;
				14'b00110000001000: oled_data = 16'b1111111111111111;
				14'b00110010001000: oled_data = 16'b1111111111111111;
				14'b00110100001000: oled_data = 16'b1111111111111111;
				14'b00110110001000: oled_data = 16'b1111111111111111;
				14'b00111000001000: oled_data = 16'b1111111111111111;
				14'b00111010001000: oled_data = 16'b1111111111111111;
				14'b00111100001000: oled_data = 16'b1111111111111111;
				14'b00111110001000: oled_data = 16'b1111111111111111;
				14'b01000000001000: oled_data = 16'b1111111111111111;
				14'b01000010001000: oled_data = 16'b1111111111111111;
				14'b01000100001000: oled_data = 16'b1111111111111111;
				14'b01000110001000: oled_data = 16'b1111111111111111;
				14'b01001000001000: oled_data = 16'b1111111111111111;
				14'b01001010001000: oled_data = 16'b1111111111111111;
				14'b01001100001000: oled_data = 16'b1111111111111111;
				14'b01001110001000: oled_data = 16'b1111111111111111;
				14'b01010000001000: oled_data = 16'b1111111111111111;
				14'b01010010001000: oled_data = 16'b1111111111111111;
				14'b01010100001000: oled_data = 16'b1111111111111111;
				14'b01010110001000: oled_data = 16'b1111111111111111;
				14'b01011000001000: oled_data = 16'b1111111111111111;
				14'b01011010001000: oled_data = 16'b1111111111111111;
				14'b01011100001000: oled_data = 16'b1111111111111111;
				14'b01011110001000: oled_data = 16'b1111111111111111;
				14'b01100000001000: oled_data = 16'b1111111111111111;
				14'b01100010001000: oled_data = 16'b1111111111111111;
				14'b01100100001000: oled_data = 16'b1111111111111111;
				14'b01100110001000: oled_data = 16'b1111111111111111;
				14'b01101000001000: oled_data = 16'b1111111111111111;
				14'b01101010001000: oled_data = 16'b1111111111111111;
				14'b01101100001000: oled_data = 16'b1111111111111111;
				14'b01101110001000: oled_data = 16'b1111111111111111;
				14'b01110000001000: oled_data = 16'b1111111111111111;
				14'b01110010001000: oled_data = 16'b1111111111111111;
				14'b01110100001000: oled_data = 16'b1111111111111111;
				14'b01110110001000: oled_data = 16'b1111111111111111;
				14'b01111000001000: oled_data = 16'b1111111111111111;
				14'b01111010001000: oled_data = 16'b1111111111111111;
				14'b01111100001000: oled_data = 16'b1111111111111111;
				14'b01111110001000: oled_data = 16'b1111111111111111;
				14'b10000000001000: oled_data = 16'b1111111111111111;
				14'b10000010001000: oled_data = 16'b1111111111111111;
				14'b10000100001000: oled_data = 16'b1111111111111111;
				14'b10000110001000: oled_data = 16'b1111111111111111;
				14'b10001000001000: oled_data = 16'b1111111111111111;
				14'b10001010001000: oled_data = 16'b1111111111111111;
				14'b10001100001000: oled_data = 16'b1111111111111111;
				14'b10001110001000: oled_data = 16'b1111111111111111;
				14'b10010000001000: oled_data = 16'b1111111111111111;
				14'b10010010001000: oled_data = 16'b1111111111111111;
				14'b10010100001000: oled_data = 16'b1111111111111111;
				14'b10010110001000: oled_data = 16'b1111111111111111;
				14'b10011000001000: oled_data = 16'b1111011111011110;
				14'b10011010001000: oled_data = 16'b1110011110011101;
				14'b10011100001000: oled_data = 16'b1101111101011100;
				14'b10011110001000: oled_data = 16'b1100111011011011;
				14'b10100000001000: oled_data = 16'b1100111011011011;
				14'b10100010001000: oled_data = 16'b1101011100111100;
				14'b10100100001000: oled_data = 16'b1101011100111100;
				14'b10100110001000: oled_data = 16'b1101111100111100;
				14'b10101000001000: oled_data = 16'b1110111110011110;
				14'b10101010001000: oled_data = 16'b1111111111111111;
				14'b10101100001000: oled_data = 16'b1111111111111111;
				14'b10101110001000: oled_data = 16'b1111111111111111;
				14'b10110000001000: oled_data = 16'b1111111111111111;
				14'b10110010001000: oled_data = 16'b1111111111111111;
				14'b10110100001000: oled_data = 16'b1111111111111111;
				14'b10110110001000: oled_data = 16'b1111111111111111;
				14'b10111000001000: oled_data = 16'b1111111111111111;
				14'b10111010001000: oled_data = 16'b1111111111111111;
				14'b10111100001000: oled_data = 16'b1111111111111111;
				14'b10111110001000: oled_data = 16'b1111111111111111;
				14'b00000000001001: oled_data = 16'b1111111111111111;
				14'b00000010001001: oled_data = 16'b1111111111111111;
				14'b00000100001001: oled_data = 16'b1111111111111111;
				14'b00000110001001: oled_data = 16'b1111111111111111;
				14'b00001000001001: oled_data = 16'b1111111111111111;
				14'b00001010001001: oled_data = 16'b1111111111111111;
				14'b00001100001001: oled_data = 16'b1111111111111111;
				14'b00001110001001: oled_data = 16'b1111111111111111;
				14'b00010000001001: oled_data = 16'b1111111111111111;
				14'b00010010001001: oled_data = 16'b1111111111111111;
				14'b00010100001001: oled_data = 16'b1111111111111111;
				14'b00010110001001: oled_data = 16'b1111111111111111;
				14'b00011000001001: oled_data = 16'b1111111111111111;
				14'b00011010001001: oled_data = 16'b1111111111111111;
				14'b00011100001001: oled_data = 16'b1111111111111111;
				14'b00011110001001: oled_data = 16'b1111111111111111;
				14'b00100000001001: oled_data = 16'b1111111111111111;
				14'b00100010001001: oled_data = 16'b1111111111111111;
				14'b00100100001001: oled_data = 16'b1111111111111111;
				14'b00100110001001: oled_data = 16'b1111111111111111;
				14'b00101000001001: oled_data = 16'b1111111111111111;
				14'b00101010001001: oled_data = 16'b1100111010011010;
				14'b00101100001001: oled_data = 16'b1101111100011011;
				14'b00101110001001: oled_data = 16'b1111111111111111;
				14'b00110000001001: oled_data = 16'b1111111111111111;
				14'b00110010001001: oled_data = 16'b1111111111111111;
				14'b00110100001001: oled_data = 16'b1111111111111111;
				14'b00110110001001: oled_data = 16'b1101011011111011;
				14'b00111000001001: oled_data = 16'b1100111010111010;
				14'b00111010001001: oled_data = 16'b1111111111111111;
				14'b00111100001001: oled_data = 16'b1111111111111111;
				14'b00111110001001: oled_data = 16'b1111111111111111;
				14'b01000000001001: oled_data = 16'b1101011010111010;
				14'b01000010001001: oled_data = 16'b1101111100011100;
				14'b01000100001001: oled_data = 16'b1111111111111111;
				14'b01000110001001: oled_data = 16'b1111111111111111;
				14'b01001000001001: oled_data = 16'b1111011111011110;
				14'b01001010001001: oled_data = 16'b1100111001111010;
				14'b01001100001001: oled_data = 16'b1111011111011110;
				14'b01001110001001: oled_data = 16'b1110111110011110;
				14'b01010000001001: oled_data = 16'b1100011001011001;
				14'b01010010001001: oled_data = 16'b1111011111011110;
				14'b01010100001001: oled_data = 16'b1111111111111111;
				14'b01010110001001: oled_data = 16'b1111111111111111;
				14'b01011000001001: oled_data = 16'b1100111010011010;
				14'b01011010001001: oled_data = 16'b1111011110111110;
				14'b01011100001001: oled_data = 16'b1111111111111111;
				14'b01011110001001: oled_data = 16'b1111111111111111;
				14'b01100000001001: oled_data = 16'b1111011111011110;
				14'b01100010001001: oled_data = 16'b1100011001011001;
				14'b01100100001001: oled_data = 16'b1110011101011101;
				14'b01100110001001: oled_data = 16'b1111111111111111;
				14'b01101000001001: oled_data = 16'b1111111111111111;
				14'b01101010001001: oled_data = 16'b1111111111111111;
				14'b01101100001001: oled_data = 16'b1111111111111111;
				14'b01101110001001: oled_data = 16'b1100111010011010;
				14'b01110000001001: oled_data = 16'b1101011011111011;
				14'b01110010001001: oled_data = 16'b1111111111111111;
				14'b01110100001001: oled_data = 16'b1110011100111100;
				14'b01110110001001: oled_data = 16'b1011010111011000;
				14'b01111000001001: oled_data = 16'b1011010111010111;
				14'b01111010001001: oled_data = 16'b1010110110110111;
				14'b01111100001001: oled_data = 16'b1101111100011100;
				14'b01111110001001: oled_data = 16'b1111111111111111;
				14'b10000000001001: oled_data = 16'b1100011001111001;
				14'b10000010001001: oled_data = 16'b1110111101111101;
				14'b10000100001001: oled_data = 16'b1111111111111111;
				14'b10000110001001: oled_data = 16'b1111111111111111;
				14'b10001000001001: oled_data = 16'b1101011011111011;
				14'b10001010001001: oled_data = 16'b1110011101011101;
				14'b10001100001001: oled_data = 16'b1111111111111111;
				14'b10001110001001: oled_data = 16'b1100111010011010;
				14'b10010000001001: oled_data = 16'b1111011110111110;
				14'b10010010001001: oled_data = 16'b1111111111111111;
				14'b10010100001001: oled_data = 16'b1111111111111111;
				14'b10010110001001: oled_data = 16'b1101011011111011;
				14'b10011000001001: oled_data = 16'b1101111100011100;
				14'b10011010001001: oled_data = 16'b1110111110011101;
				14'b10011100001001: oled_data = 16'b1110011101111101;
				14'b10011110001001: oled_data = 16'b1100111011111011;
				14'b10100000001001: oled_data = 16'b1100111011011011;
				14'b10100010001001: oled_data = 16'b1101011100011011;
				14'b10100100001001: oled_data = 16'b1101111100111100;
				14'b10100110001001: oled_data = 16'b1101011100111100;
				14'b10101000001001: oled_data = 16'b1110011101111101;
				14'b10101010001001: oled_data = 16'b1111011111011110;
				14'b10101100001001: oled_data = 16'b1111111111111111;
				14'b10101110001001: oled_data = 16'b1111111111111111;
				14'b10110000001001: oled_data = 16'b1111111111111111;
				14'b10110010001001: oled_data = 16'b1111111111111111;
				14'b10110100001001: oled_data = 16'b1111111111111111;
				14'b10110110001001: oled_data = 16'b1111111111111111;
				14'b10111000001001: oled_data = 16'b1111111111111111;
				14'b10111010001001: oled_data = 16'b1111111111111111;
				14'b10111100001001: oled_data = 16'b1111111111111111;
				14'b10111110001001: oled_data = 16'b1111111111111111;
				14'b00000000001010: oled_data = 16'b1111111111111111;
				14'b00000010001010: oled_data = 16'b1111111111111111;
				14'b00000100001010: oled_data = 16'b1111111111111111;
				14'b00000110001010: oled_data = 16'b1111111111111111;
				14'b00001000001010: oled_data = 16'b1111111111111111;
				14'b00001010001010: oled_data = 16'b1111111111111111;
				14'b00001100001010: oled_data = 16'b1111111111111111;
				14'b00001110001010: oled_data = 16'b1111111111111111;
				14'b00010000001010: oled_data = 16'b1111111111111111;
				14'b00010010001010: oled_data = 16'b1111111111111111;
				14'b00010100001010: oled_data = 16'b1111111111111111;
				14'b00010110001010: oled_data = 16'b1111111111111111;
				14'b00011000001010: oled_data = 16'b1111111111111111;
				14'b00011010001010: oled_data = 16'b1111111111111111;
				14'b00011100001010: oled_data = 16'b1111111111111111;
				14'b00011110001010: oled_data = 16'b1111111111111111;
				14'b00100000001010: oled_data = 16'b1111111111111111;
				14'b00100010001010: oled_data = 16'b1111111111111111;
				14'b00100100001010: oled_data = 16'b1111111111111111;
				14'b00100110001010: oled_data = 16'b1111111111111111;
				14'b00101000001010: oled_data = 16'b1111111111111111;
				14'b00101010001010: oled_data = 16'b0110001101101111;
				14'b00101100001010: oled_data = 16'b0110001110010000;
				14'b00101110001010: oled_data = 16'b1111011111011110;
				14'b00110000001010: oled_data = 16'b1111111111111111;
				14'b00110010001010: oled_data = 16'b1111111111111111;
				14'b00110100001010: oled_data = 16'b1111011110111110;
				14'b00110110001010: oled_data = 16'b0101101101001111;
				14'b00111000001010: oled_data = 16'b0110101111010001;
				14'b00111010001010: oled_data = 16'b1111111111111111;
				14'b00111100001010: oled_data = 16'b1111111111111111;
				14'b00111110001010: oled_data = 16'b1111011111011110;
				14'b01000000001010: oled_data = 16'b0101101101101111;
				14'b01000010001010: oled_data = 16'b0111110001010010;
				14'b01000100001010: oled_data = 16'b1111111111111111;
				14'b01000110001010: oled_data = 16'b1111111111111111;
				14'b01001000001010: oled_data = 16'b1110111110011101;
				14'b01001010001010: oled_data = 16'b0110101110110000;
				14'b01001100001010: oled_data = 16'b1111011110111110;
				14'b01001110001010: oled_data = 16'b1101011011011011;
				14'b01010000001010: oled_data = 16'b0011101001001100;
				14'b01010010001010: oled_data = 16'b1010110110010111;
				14'b01010100001010: oled_data = 16'b1111111111111111;
				14'b01010110001010: oled_data = 16'b1111011111011110;
				14'b01011000001010: oled_data = 16'b0110101111010001;
				14'b01011010001010: oled_data = 16'b1101111100011100;
				14'b01011100001010: oled_data = 16'b1111111111111111;
				14'b01011110001010: oled_data = 16'b1111111111111111;
				14'b01100000001010: oled_data = 16'b1110111110011101;
				14'b01100010001010: oled_data = 16'b0100101011001101;
				14'b01100100001010: oled_data = 16'b1000010001110011;
				14'b01100110001010: oled_data = 16'b1111111111111111;
				14'b01101000001010: oled_data = 16'b1111111111111111;
				14'b01101010001010: oled_data = 16'b1111111111111111;
				14'b01101100001010: oled_data = 16'b1110011101011101;
				14'b01101110001010: oled_data = 16'b0100001010101101;
				14'b01110000001010: oled_data = 16'b1000110010110100;
				14'b01110010001010: oled_data = 16'b1111111111111111;
				14'b01110100001010: oled_data = 16'b1010010101010110;
				14'b01110110001010: oled_data = 16'b0110101111010001;
				14'b01111000001010: oled_data = 16'b1001110100110101;
				14'b01111010001010: oled_data = 16'b1001110100010101;
				14'b01111100001010: oled_data = 16'b1101011011011011;
				14'b01111110001010: oled_data = 16'b1111011110111110;
				14'b10000000001010: oled_data = 16'b0100101011101101;
				14'b10000010001010: oled_data = 16'b0111110001010010;
				14'b10000100001010: oled_data = 16'b1111111111111111;
				14'b10000110001010: oled_data = 16'b1111111111111111;
				14'b10001000001010: oled_data = 16'b1000110010010011;
				14'b10001010001010: oled_data = 16'b1011010111111000;
				14'b10001100001010: oled_data = 16'b1111111111111111;
				14'b10001110001010: oled_data = 16'b0110101110110000;
				14'b10010000001010: oled_data = 16'b1110011101011100;
				14'b10010010001010: oled_data = 16'b1111111111111111;
				14'b10010100001010: oled_data = 16'b1111111111111111;
				14'b10010110001010: oled_data = 16'b1001010011110101;
				14'b10011000001010: oled_data = 16'b1010010110010110;
				14'b10011010001010: oled_data = 16'b1111011111011110;
				14'b10011100001010: oled_data = 16'b1110011110011101;
				14'b10011110001010: oled_data = 16'b1101011100011011;
				14'b10100000001010: oled_data = 16'b1100111011011010;
				14'b10100010001010: oled_data = 16'b1100111011111011;
				14'b10100100001010: oled_data = 16'b1101111100111100;
				14'b10100110001010: oled_data = 16'b1101111100111100;
				14'b10101000001010: oled_data = 16'b1101111101011100;
				14'b10101010001010: oled_data = 16'b1110111110011110;
				14'b10101100001010: oled_data = 16'b1111111111111111;
				14'b10101110001010: oled_data = 16'b1111111111111111;
				14'b10110000001010: oled_data = 16'b1111111111111111;
				14'b10110010001010: oled_data = 16'b1111111111111111;
				14'b10110100001010: oled_data = 16'b1111111111111111;
				14'b10110110001010: oled_data = 16'b1111111111111111;
				14'b10111000001010: oled_data = 16'b1111111111111111;
				14'b10111010001010: oled_data = 16'b1111111111111111;
				14'b10111100001010: oled_data = 16'b1111111111111111;
				14'b10111110001010: oled_data = 16'b1111111111111111;
				14'b00000000001011: oled_data = 16'b1111111111111111;
				14'b00000010001011: oled_data = 16'b1111111111111111;
				14'b00000100001011: oled_data = 16'b1111111111111111;
				14'b00000110001011: oled_data = 16'b1111111111111111;
				14'b00001000001011: oled_data = 16'b1111111111111111;
				14'b00001010001011: oled_data = 16'b1111111111111111;
				14'b00001100001011: oled_data = 16'b1111111111111111;
				14'b00001110001011: oled_data = 16'b1111111111111111;
				14'b00010000001011: oled_data = 16'b1111111111111111;
				14'b00010010001011: oled_data = 16'b1111111111111111;
				14'b00010100001011: oled_data = 16'b1111111111111111;
				14'b00010110001011: oled_data = 16'b1111111111111111;
				14'b00011000001011: oled_data = 16'b1111111111111111;
				14'b00011010001011: oled_data = 16'b1111111111111111;
				14'b00011100001011: oled_data = 16'b1111111111111111;
				14'b00011110001011: oled_data = 16'b1111111111111111;
				14'b00100000001011: oled_data = 16'b1111111111111111;
				14'b00100010001011: oled_data = 16'b1111111111111111;
				14'b00100100001011: oled_data = 16'b1111111111111111;
				14'b00100110001011: oled_data = 16'b1111111111111111;
				14'b00101000001011: oled_data = 16'b1111011111011110;
				14'b00101010001011: oled_data = 16'b0111010000010001;
				14'b00101100001011: oled_data = 16'b0101101101101111;
				14'b00101110001011: oled_data = 16'b1100111010011010;
				14'b00110000001011: oled_data = 16'b1111111111111111;
				14'b00110010001011: oled_data = 16'b1111111111111111;
				14'b00110100001011: oled_data = 16'b1011111000111001;
				14'b00110110001011: oled_data = 16'b0110001110010000;
				14'b00111000001011: oled_data = 16'b0111110001010010;
				14'b00111010001011: oled_data = 16'b1111111111111111;
				14'b00111100001011: oled_data = 16'b1111111111111111;
				14'b00111110001011: oled_data = 16'b1100111010011010;
				14'b01000000001011: oled_data = 16'b0111110001010010;
				14'b01000010001011: oled_data = 16'b0111010000010001;
				14'b01000100001011: oled_data = 16'b1110011100111100;
				14'b01000110001011: oled_data = 16'b1111111111111111;
				14'b01001000001011: oled_data = 16'b1110111110011101;
				14'b01001010001011: oled_data = 16'b0110101111010001;
				14'b01001100001011: oled_data = 16'b1111011110111110;
				14'b01001110001011: oled_data = 16'b1101011010111010;
				14'b01010000001011: oled_data = 16'b0110001110010000;
				14'b01010010001011: oled_data = 16'b0110101110110000;
				14'b01010100001011: oled_data = 16'b1110011101011101;
				14'b01010110001011: oled_data = 16'b1111111111111111;
				14'b01011000001011: oled_data = 16'b0111001111110001;
				14'b01011010001011: oled_data = 16'b1101111100011100;
				14'b01011100001011: oled_data = 16'b1111111111111111;
				14'b01011110001011: oled_data = 16'b1111111111111111;
				14'b01100000001011: oled_data = 16'b1110111101111101;
				14'b01100010001011: oled_data = 16'b0110001110110000;
				14'b01100100001011: oled_data = 16'b0110001110010000;
				14'b01100110001011: oled_data = 16'b1101111100111100;
				14'b01101000001011: oled_data = 16'b1111111111111111;
				14'b01101010001011: oled_data = 16'b1111111111111111;
				14'b01101100001011: oled_data = 16'b1010010101110110;
				14'b01101110001011: oled_data = 16'b0110001110010000;
				14'b01110000001011: oled_data = 16'b1001010011110100;
				14'b01110010001011: oled_data = 16'b1111111111111111;
				14'b01110100001011: oled_data = 16'b1001110100110101;
				14'b01110110001011: oled_data = 16'b1010110110010111;
				14'b01111000001011: oled_data = 16'b1111111111111111;
				14'b01111010001011: oled_data = 16'b1111111111111111;
				14'b01111100001011: oled_data = 16'b1111111111111111;
				14'b01111110001011: oled_data = 16'b1110111110011101;
				14'b10000000001011: oled_data = 16'b0110101111010000;
				14'b10000010001011: oled_data = 16'b0110001110010000;
				14'b10000100001011: oled_data = 16'b1100011001111010;
				14'b10000110001011: oled_data = 16'b1111111111111111;
				14'b10001000001011: oled_data = 16'b1000110010110100;
				14'b10001010001011: oled_data = 16'b1011011000011000;
				14'b10001100001011: oled_data = 16'b1111111111111111;
				14'b10001110001011: oled_data = 16'b0110101111010001;
				14'b10010000001011: oled_data = 16'b1110011101011100;
				14'b10010010001011: oled_data = 16'b1111111111111111;
				14'b10010100001011: oled_data = 16'b1111111111111111;
				14'b10010110001011: oled_data = 16'b1001010100010101;
				14'b10011000001011: oled_data = 16'b1010110110010111;
				14'b10011010001011: oled_data = 16'b1111111111111111;
				14'b10011100001011: oled_data = 16'b1110111110011101;
				14'b10011110001011: oled_data = 16'b1110011101011100;
				14'b10100000001011: oled_data = 16'b1100111011011010;
				14'b10100010001011: oled_data = 16'b1100111011011010;
				14'b10100100001011: oled_data = 16'b1101011100011011;
				14'b10100110001011: oled_data = 16'b1101111100111100;
				14'b10101000001011: oled_data = 16'b1101111100111100;
				14'b10101010001011: oled_data = 16'b1110011101111101;
				14'b10101100001011: oled_data = 16'b1111011111011110;
				14'b10101110001011: oled_data = 16'b1111111111111111;
				14'b10110000001011: oled_data = 16'b1111111111111111;
				14'b10110010001011: oled_data = 16'b1111111111111111;
				14'b10110100001011: oled_data = 16'b1111111111111111;
				14'b10110110001011: oled_data = 16'b1111111111111111;
				14'b10111000001011: oled_data = 16'b1111111111111111;
				14'b10111010001011: oled_data = 16'b1111111111111111;
				14'b10111100001011: oled_data = 16'b1111111111111111;
				14'b10111110001011: oled_data = 16'b1111111111111111;
				14'b00000000001100: oled_data = 16'b1111111111111111;
				14'b00000010001100: oled_data = 16'b1111111111111111;
				14'b00000100001100: oled_data = 16'b1111111111111111;
				14'b00000110001100: oled_data = 16'b1111111111111111;
				14'b00001000001100: oled_data = 16'b1111111111111111;
				14'b00001010001100: oled_data = 16'b1111111111111111;
				14'b00001100001100: oled_data = 16'b1111111111111111;
				14'b00001110001100: oled_data = 16'b1111111111111111;
				14'b00010000001100: oled_data = 16'b1111111111111111;
				14'b00010010001100: oled_data = 16'b1111111111111111;
				14'b00010100001100: oled_data = 16'b1111111111111111;
				14'b00010110001100: oled_data = 16'b1111111111111111;
				14'b00011000001100: oled_data = 16'b1111111111111111;
				14'b00011010001100: oled_data = 16'b1111111111111111;
				14'b00011100001100: oled_data = 16'b1111111111111111;
				14'b00011110001100: oled_data = 16'b1111111111111111;
				14'b00100000001100: oled_data = 16'b1111111111111111;
				14'b00100010001100: oled_data = 16'b1111111111111111;
				14'b00100100001100: oled_data = 16'b1111111111111111;
				14'b00100110001100: oled_data = 16'b1111111111111111;
				14'b00101000001100: oled_data = 16'b1111011111011110;
				14'b00101010001100: oled_data = 16'b0111010000010010;
				14'b00101100001100: oled_data = 16'b1010010101010110;
				14'b00101110001100: oled_data = 16'b1000010001110011;
				14'b00110000001100: oled_data = 16'b1111111111111111;
				14'b00110010001100: oled_data = 16'b1111011111011110;
				14'b00110100001100: oled_data = 16'b0111110001010010;
				14'b00110110001100: oled_data = 16'b1010110110010111;
				14'b00111000001100: oled_data = 16'b0111110000110010;
				14'b00111010001100: oled_data = 16'b1111111111111111;
				14'b00111100001100: oled_data = 16'b1111111111111111;
				14'b00111110001100: oled_data = 16'b1000110010110100;
				14'b01000000001100: oled_data = 16'b1100011001111001;
				14'b01000010001100: oled_data = 16'b1010010101010110;
				14'b01000100001100: oled_data = 16'b1010010110010110;
				14'b01000110001100: oled_data = 16'b1111111111111111;
				14'b01001000001100: oled_data = 16'b1110111110011101;
				14'b01001010001100: oled_data = 16'b0110101111010001;
				14'b01001100001100: oled_data = 16'b1111011110111110;
				14'b01001110001100: oled_data = 16'b1100111010111010;
				14'b01010000001100: oled_data = 16'b1000010001110011;
				14'b01010010001100: oled_data = 16'b1010010101110110;
				14'b01010100001100: oled_data = 16'b1000110011010100;
				14'b01010110001100: oled_data = 16'b1111111111111111;
				14'b01011000001100: oled_data = 16'b0111001111110001;
				14'b01011010001100: oled_data = 16'b1101111100011100;
				14'b01011100001100: oled_data = 16'b1111111111111111;
				14'b01011110001100: oled_data = 16'b1111111111111111;
				14'b01100000001100: oled_data = 16'b1110011101111101;
				14'b01100010001100: oled_data = 16'b0111010000010001;
				14'b01100100001100: oled_data = 16'b1001010100010101;
				14'b01100110001100: oled_data = 16'b1001110100110101;
				14'b01101000001100: oled_data = 16'b1111111111111111;
				14'b01101010001100: oled_data = 16'b1110111110011110;
				14'b01101100001100: oled_data = 16'b0111010000010001;
				14'b01101110001100: oled_data = 16'b1010010101110110;
				14'b01110000001100: oled_data = 16'b1000110011010100;
				14'b01110010001100: oled_data = 16'b1111111111111111;
				14'b01110100001100: oled_data = 16'b1010010101010110;
				14'b01110110001100: oled_data = 16'b1000010001110011;
				14'b01111000001100: oled_data = 16'b1011111000011001;
				14'b01111010001100: oled_data = 16'b1100011001011001;
				14'b01111100001100: oled_data = 16'b1111011110111110;
				14'b01111110001100: oled_data = 16'b1110111110011101;
				14'b10000000001100: oled_data = 16'b0111001111110001;
				14'b10000010001100: oled_data = 16'b1011111000111001;
				14'b10000100001100: oled_data = 16'b0110101111110001;
				14'b10000110001100: oled_data = 16'b1111011111011110;
				14'b10001000001100: oled_data = 16'b1000110010110100;
				14'b10001010001100: oled_data = 16'b1011011000011000;
				14'b10001100001100: oled_data = 16'b1111111111111111;
				14'b10001110001100: oled_data = 16'b0110101111010001;
				14'b10010000001100: oled_data = 16'b1110011101011100;
				14'b10010010001100: oled_data = 16'b1111111111111111;
				14'b10010100001100: oled_data = 16'b1111111111111111;
				14'b10010110001100: oled_data = 16'b1001010100010101;
				14'b10011000001100: oled_data = 16'b1010110110010111;
				14'b10011010001100: oled_data = 16'b1111111111111111;
				14'b10011100001100: oled_data = 16'b1110111110111101;
				14'b10011110001100: oled_data = 16'b1110011110011101;
				14'b10100000001100: oled_data = 16'b1101011100011011;
				14'b10100010001100: oled_data = 16'b1100111011111010;
				14'b10100100001100: oled_data = 16'b1101011011111011;
				14'b10100110001100: oled_data = 16'b1101111100111100;
				14'b10101000001100: oled_data = 16'b1101111100111100;
				14'b10101010001100: oled_data = 16'b1101111100111100;
				14'b10101100001100: oled_data = 16'b1110111110011101;
				14'b10101110001100: oled_data = 16'b1111011111111111;
				14'b10110000001100: oled_data = 16'b1111111111111111;
				14'b10110010001100: oled_data = 16'b1111111111111111;
				14'b10110100001100: oled_data = 16'b1111111111111111;
				14'b10110110001100: oled_data = 16'b1111111111111111;
				14'b10111000001100: oled_data = 16'b1111111111111111;
				14'b10111010001100: oled_data = 16'b1111111111111111;
				14'b10111100001100: oled_data = 16'b1111111111111111;
				14'b10111110001100: oled_data = 16'b1111111111111111;
				14'b00000000001101: oled_data = 16'b1111111111111111;
				14'b00000010001101: oled_data = 16'b1111111111111111;
				14'b00000100001101: oled_data = 16'b1111111111111111;
				14'b00000110001101: oled_data = 16'b1111111111111111;
				14'b00001000001101: oled_data = 16'b1111111111111111;
				14'b00001010001101: oled_data = 16'b1111111111111111;
				14'b00001100001101: oled_data = 16'b1111111111111111;
				14'b00001110001101: oled_data = 16'b1111111111111111;
				14'b00010000001101: oled_data = 16'b1111111111111111;
				14'b00010010001101: oled_data = 16'b1111111111111111;
				14'b00010100001101: oled_data = 16'b1111111111111111;
				14'b00010110001101: oled_data = 16'b1111111111111111;
				14'b00011000001101: oled_data = 16'b1111111111111111;
				14'b00011010001101: oled_data = 16'b1111111111111111;
				14'b00011100001101: oled_data = 16'b1111111111111111;
				14'b00011110001101: oled_data = 16'b1111111111111111;
				14'b00100000001101: oled_data = 16'b1111111111111111;
				14'b00100010001101: oled_data = 16'b1111111111111111;
				14'b00100100001101: oled_data = 16'b1111111111111111;
				14'b00100110001101: oled_data = 16'b1111111111111111;
				14'b00101000001101: oled_data = 16'b1111011111011110;
				14'b00101010001101: oled_data = 16'b0111001111110001;
				14'b00101100001101: oled_data = 16'b1101011011111011;
				14'b00101110001101: oled_data = 16'b0110101111010001;
				14'b00110000001101: oled_data = 16'b1110011100111100;
				14'b00110010001101: oled_data = 16'b1101011011011011;
				14'b00110100001101: oled_data = 16'b0111110001010010;
				14'b00110110001101: oled_data = 16'b1101011011011011;
				14'b00111000001101: oled_data = 16'b0111010000010010;
				14'b00111010001101: oled_data = 16'b1111111111111111;
				14'b00111100001101: oled_data = 16'b1110111110011101;
				14'b00111110001101: oled_data = 16'b0110101111110001;
				14'b01000000001101: oled_data = 16'b1110111110011101;
				14'b01000010001101: oled_data = 16'b1101011011011011;
				14'b01000100001101: oled_data = 16'b0111010000010001;
				14'b01000110001101: oled_data = 16'b1111011111011110;
				14'b01001000001101: oled_data = 16'b1110111110011101;
				14'b01001010001101: oled_data = 16'b0110101111010001;
				14'b01001100001101: oled_data = 16'b1111011110111110;
				14'b01001110001101: oled_data = 16'b1100111010111010;
				14'b01010000001101: oled_data = 16'b0111110001010010;
				14'b01010010001101: oled_data = 16'b1111011110111110;
				14'b01010100001101: oled_data = 16'b0110101110110000;
				14'b01010110001101: oled_data = 16'b1101011011011011;
				14'b01011000001101: oled_data = 16'b0111010000010001;
				14'b01011010001101: oled_data = 16'b1101111100011100;
				14'b01011100001101: oled_data = 16'b1111111111111111;
				14'b01011110001101: oled_data = 16'b1111111111111111;
				14'b01100000001101: oled_data = 16'b1110011101111101;
				14'b01100010001101: oled_data = 16'b0110101111110001;
				14'b01100100001101: oled_data = 16'b1101111011111011;
				14'b01100110001101: oled_data = 16'b0110101111010000;
				14'b01101000001101: oled_data = 16'b1111011110111110;
				14'b01101010001101: oled_data = 16'b1011010111111000;
				14'b01101100001101: oled_data = 16'b1001010100010101;
				14'b01101110001101: oled_data = 16'b1011111000111001;
				14'b01110000001101: oled_data = 16'b1000110010110100;
				14'b01110010001101: oled_data = 16'b1111111111111111;
				14'b01110100001101: oled_data = 16'b1010010101010110;
				14'b01110110001101: oled_data = 16'b0110101111010000;
				14'b01111000001101: oled_data = 16'b1001010100010101;
				14'b01111010001101: oled_data = 16'b1001110100110101;
				14'b01111100001101: oled_data = 16'b1110111110011110;
				14'b01111110001101: oled_data = 16'b1110111110011101;
				14'b10000000001101: oled_data = 16'b0110101111010001;
				14'b10000010001101: oled_data = 16'b1111011110111110;
				14'b10000100001101: oled_data = 16'b1000010001110011;
				14'b10000110001101: oled_data = 16'b1011010111111000;
				14'b10001000001101: oled_data = 16'b1001010011110100;
				14'b10001010001101: oled_data = 16'b1011011000011000;
				14'b10001100001101: oled_data = 16'b1111111111111111;
				14'b10001110001101: oled_data = 16'b0110101111010001;
				14'b10010000001101: oled_data = 16'b1110011101011100;
				14'b10010010001101: oled_data = 16'b1111111111111111;
				14'b10010100001101: oled_data = 16'b1111111111111111;
				14'b10010110001101: oled_data = 16'b1001110100010101;
				14'b10011000001101: oled_data = 16'b1010110110010111;
				14'b10011010001101: oled_data = 16'b1111111111111111;
				14'b10011100001101: oled_data = 16'b1111011111011110;
				14'b10011110001101: oled_data = 16'b1110111110011101;
				14'b10100000001101: oled_data = 16'b1101111101111100;
				14'b10100010001101: oled_data = 16'b1100111011111010;
				14'b10100100001101: oled_data = 16'b1100111100011010;
				14'b10100110001101: oled_data = 16'b1101011100111011;
				14'b10101000001101: oled_data = 16'b1101111100111100;
				14'b10101010001101: oled_data = 16'b1101111100111100;
				14'b10101100001101: oled_data = 16'b1110011101111100;
				14'b10101110001101: oled_data = 16'b1111011110111110;
				14'b10110000001101: oled_data = 16'b1111111111111111;
				14'b10110010001101: oled_data = 16'b1111111111111111;
				14'b10110100001101: oled_data = 16'b1111111111111111;
				14'b10110110001101: oled_data = 16'b1111111111111111;
				14'b10111000001101: oled_data = 16'b1111111111111111;
				14'b10111010001101: oled_data = 16'b1111111111111111;
				14'b10111100001101: oled_data = 16'b1111111111111111;
				14'b10111110001101: oled_data = 16'b1111111111111111;
				14'b00000000001110: oled_data = 16'b1111111111111111;
				14'b00000010001110: oled_data = 16'b1111111111111111;
				14'b00000100001110: oled_data = 16'b1111111111111111;
				14'b00000110001110: oled_data = 16'b1111111111111111;
				14'b00001000001110: oled_data = 16'b1111111111111111;
				14'b00001010001110: oled_data = 16'b1111111111111111;
				14'b00001100001110: oled_data = 16'b1111111111111111;
				14'b00001110001110: oled_data = 16'b1111111111111111;
				14'b00010000001110: oled_data = 16'b1111111111111111;
				14'b00010010001110: oled_data = 16'b1111111111111111;
				14'b00010100001110: oled_data = 16'b1111111111111111;
				14'b00010110001110: oled_data = 16'b1111111111111111;
				14'b00011000001110: oled_data = 16'b1111111111111111;
				14'b00011010001110: oled_data = 16'b1111111111111111;
				14'b00011100001110: oled_data = 16'b1111111111111111;
				14'b00011110001110: oled_data = 16'b1111111111111111;
				14'b00100000001110: oled_data = 16'b1111111111111111;
				14'b00100010001110: oled_data = 16'b1111111111111111;
				14'b00100100001110: oled_data = 16'b1111111111111111;
				14'b00100110001110: oled_data = 16'b1111111111111111;
				14'b00101000001110: oled_data = 16'b1111011111011110;
				14'b00101010001110: oled_data = 16'b0110101111110001;
				14'b00101100001110: oled_data = 16'b1110011101011101;
				14'b00101110001110: oled_data = 16'b1010010101010110;
				14'b00110000001110: oled_data = 16'b1001110100110101;
				14'b00110010001110: oled_data = 16'b1000110011010100;
				14'b00110100001110: oled_data = 16'b1100011001011001;
				14'b00110110001110: oled_data = 16'b1101011011111011;
				14'b00111000001110: oled_data = 16'b0111010000010010;
				14'b00111010001110: oled_data = 16'b1111111111111111;
				14'b00111100001110: oled_data = 16'b1011111000111001;
				14'b00111110001110: oled_data = 16'b0101001100001110;
				14'b01000000001110: oled_data = 16'b0111110001010010;
				14'b01000010001110: oled_data = 16'b0111110000110010;
				14'b01000100001110: oled_data = 16'b0101001100001110;
				14'b01000110001110: oled_data = 16'b1101011011111011;
				14'b01001000001110: oled_data = 16'b1111011110111110;
				14'b01001010001110: oled_data = 16'b0110101111010001;
				14'b01001100001110: oled_data = 16'b1111011110111110;
				14'b01001110001110: oled_data = 16'b1100111010111010;
				14'b01010000001110: oled_data = 16'b0111110000110010;
				14'b01010010001110: oled_data = 16'b1111111111111111;
				14'b01010100001110: oled_data = 16'b1011010111111000;
				14'b01010110001110: oled_data = 16'b0111110000110010;
				14'b01011000001110: oled_data = 16'b0111010000010001;
				14'b01011010001110: oled_data = 16'b1101111100011100;
				14'b01011100001110: oled_data = 16'b1111111111111111;
				14'b01011110001110: oled_data = 16'b1111111111111111;
				14'b01100000001110: oled_data = 16'b1110011101111101;
				14'b01100010001110: oled_data = 16'b0110101111010001;
				14'b01100100001110: oled_data = 16'b1111011111011110;
				14'b01100110001110: oled_data = 16'b1000010010010011;
				14'b01101000001110: oled_data = 16'b1011010111010111;
				14'b01101010001110: oled_data = 16'b0111110001010010;
				14'b01101100001110: oled_data = 16'b1101111100011100;
				14'b01101110001110: oled_data = 16'b1011111000011000;
				14'b01110000001110: oled_data = 16'b1000110010110100;
				14'b01110010001110: oled_data = 16'b1111111111111111;
				14'b01110100001110: oled_data = 16'b1001110101010110;
				14'b01110110001110: oled_data = 16'b1010010110010110;
				14'b01111000001110: oled_data = 16'b1111111111111111;
				14'b01111010001110: oled_data = 16'b1111111111111111;
				14'b01111100001110: oled_data = 16'b1111111111111111;
				14'b01111110001110: oled_data = 16'b1110111110011101;
				14'b10000000001110: oled_data = 16'b0110101111010001;
				14'b10000010001110: oled_data = 16'b1111011110111110;
				14'b10000100001110: oled_data = 16'b1101111100011100;
				14'b10000110001110: oled_data = 16'b0110101111010001;
				14'b10001000001110: oled_data = 16'b0111110001010010;
				14'b10001010001110: oled_data = 16'b1011111000011000;
				14'b10001100001110: oled_data = 16'b1111111111111111;
				14'b10001110001110: oled_data = 16'b0110101111010001;
				14'b10010000001110: oled_data = 16'b1110011101011100;
				14'b10010010001110: oled_data = 16'b1111111111111111;
				14'b10010100001110: oled_data = 16'b1111111111111111;
				14'b10010110001110: oled_data = 16'b1001010011110101;
				14'b10011000001110: oled_data = 16'b1010110110110111;
				14'b10011010001110: oled_data = 16'b1111111111111111;
				14'b10011100001110: oled_data = 16'b1111111111111111;
				14'b10011110001110: oled_data = 16'b1110111110111101;
				14'b10100000001110: oled_data = 16'b1110011110011101;
				14'b10100010001110: oled_data = 16'b1101011100111011;
				14'b10100100001110: oled_data = 16'b1100111100011010;
				14'b10100110001110: oled_data = 16'b1101011100011010;
				14'b10101000001110: oled_data = 16'b1101111101011100;
				14'b10101010001110: oled_data = 16'b1101111101011100;
				14'b10101100001110: oled_data = 16'b1101111101011100;
				14'b10101110001110: oled_data = 16'b1110011110011101;
				14'b10110000001110: oled_data = 16'b1111011111011110;
				14'b10110010001110: oled_data = 16'b1111111111111111;
				14'b10110100001110: oled_data = 16'b1111111111111111;
				14'b10110110001110: oled_data = 16'b1111111111111111;
				14'b10111000001110: oled_data = 16'b1111111111111111;
				14'b10111010001110: oled_data = 16'b1111111111111111;
				14'b10111100001110: oled_data = 16'b1111111111111111;
				14'b10111110001110: oled_data = 16'b1111111111111111;
				14'b00000000001111: oled_data = 16'b1111111111111111;
				14'b00000010001111: oled_data = 16'b1111111111111111;
				14'b00000100001111: oled_data = 16'b1111111111111111;
				14'b00000110001111: oled_data = 16'b1111111111111111;
				14'b00001000001111: oled_data = 16'b1111111111111111;
				14'b00001010001111: oled_data = 16'b1111111111111111;
				14'b00001100001111: oled_data = 16'b1111111111111111;
				14'b00001110001111: oled_data = 16'b1111111111111111;
				14'b00010000001111: oled_data = 16'b1111111111111111;
				14'b00010010001111: oled_data = 16'b1111111111111111;
				14'b00010100001111: oled_data = 16'b1111111111111111;
				14'b00010110001111: oled_data = 16'b1111111111111111;
				14'b00011000001111: oled_data = 16'b1111111111111111;
				14'b00011010001111: oled_data = 16'b1111111111111111;
				14'b00011100001111: oled_data = 16'b1111111111111111;
				14'b00011110001111: oled_data = 16'b1111111111111111;
				14'b00100000001111: oled_data = 16'b1111111111111111;
				14'b00100010001111: oled_data = 16'b1111111111111111;
				14'b00100100001111: oled_data = 16'b1111111111111111;
				14'b00100110001111: oled_data = 16'b1111111111111111;
				14'b00101000001111: oled_data = 16'b1111011111011110;
				14'b00101010001111: oled_data = 16'b0110101111010001;
				14'b00101100001111: oled_data = 16'b1101111100111100;
				14'b00101110001111: oled_data = 16'b1110011101011101;
				14'b00110000001111: oled_data = 16'b0101001100101110;
				14'b00110010001111: oled_data = 16'b0110101111010001;
				14'b00110100001111: oled_data = 16'b1111011111011110;
				14'b00110110001111: oled_data = 16'b1101011011011011;
				14'b00111000001111: oled_data = 16'b0111010000010001;
				14'b00111010001111: oled_data = 16'b1111111111111111;
				14'b00111100001111: oled_data = 16'b0111110000110010;
				14'b00111110001111: oled_data = 16'b1011111000011000;
				14'b01000000001111: oled_data = 16'b1110111110011101;
				14'b01000010001111: oled_data = 16'b1110111110011101;
				14'b01000100001111: oled_data = 16'b1001110101010110;
				14'b01000110001111: oled_data = 16'b1001010011110100;
				14'b01001000001111: oled_data = 16'b1111011110111110;
				14'b01001010001111: oled_data = 16'b0110101110110000;
				14'b01001100001111: oled_data = 16'b1111011110111110;
				14'b01001110001111: oled_data = 16'b1100111010011010;
				14'b01010000001111: oled_data = 16'b0111010000110010;
				14'b01010010001111: oled_data = 16'b1111111111111111;
				14'b01010100001111: oled_data = 16'b1111011111011110;
				14'b01010110001111: oled_data = 16'b0111010000010001;
				14'b01011000001111: oled_data = 16'b0100001010101101;
				14'b01011010001111: oled_data = 16'b1101111100111100;
				14'b01011100001111: oled_data = 16'b1111111111111111;
				14'b01011110001111: oled_data = 16'b1111111111111111;
				14'b01100000001111: oled_data = 16'b1110011101111101;
				14'b01100010001111: oled_data = 16'b0110101110110000;
				14'b01100100001111: oled_data = 16'b1111011111011110;
				14'b01100110001111: oled_data = 16'b1100111010111010;
				14'b01101000001111: oled_data = 16'b0100101011101101;
				14'b01101010001111: oled_data = 16'b1000010001110011;
				14'b01101100001111: oled_data = 16'b1111111111111111;
				14'b01101110001111: oled_data = 16'b1011010111111000;
				14'b01110000001111: oled_data = 16'b1000110010110011;
				14'b01110010001111: oled_data = 16'b1111111111111111;
				14'b01110100001111: oled_data = 16'b1001110100110101;
				14'b01110110001111: oled_data = 16'b1001110100110101;
				14'b01111000001111: oled_data = 16'b1110111110011101;
				14'b01111010001111: oled_data = 16'b1110111110011101;
				14'b01111100001111: oled_data = 16'b1111011111011110;
				14'b01111110001111: oled_data = 16'b1110111110011101;
				14'b10000000001111: oled_data = 16'b0110101110110000;
				14'b10000010001111: oled_data = 16'b1110111110011101;
				14'b10000100001111: oled_data = 16'b1111111111111111;
				14'b10000110001111: oled_data = 16'b1001110100110101;
				14'b10001000001111: oled_data = 16'b0011101001101100;
				14'b10001010001111: oled_data = 16'b1011111000111001;
				14'b10001100001111: oled_data = 16'b1111111111111111;
				14'b10001110001111: oled_data = 16'b1000010001110011;
				14'b10010000001111: oled_data = 16'b1001110101010110;
				14'b10010010001111: oled_data = 16'b1111011110111110;
				14'b10010100001111: oled_data = 16'b1110011100111100;
				14'b10010110001111: oled_data = 16'b0110101110110000;
				14'b10011000001111: oled_data = 16'b1101011011011011;
				14'b10011010001111: oled_data = 16'b1111111111111111;
				14'b10011100001111: oled_data = 16'b1111111111111111;
				14'b10011110001111: oled_data = 16'b1111011111011110;
				14'b10100000001111: oled_data = 16'b1110111110011101;
				14'b10100010001111: oled_data = 16'b1110011101111100;
				14'b10100100001111: oled_data = 16'b1100111011111010;
				14'b10100110001111: oled_data = 16'b1100111100011010;
				14'b10101000001111: oled_data = 16'b1101011100111011;
				14'b10101010001111: oled_data = 16'b1101111101011011;
				14'b10101100001111: oled_data = 16'b1101111101011011;
				14'b10101110001111: oled_data = 16'b1101111101011100;
				14'b10110000001111: oled_data = 16'b1110111110011101;
				14'b10110010001111: oled_data = 16'b1111011111011110;
				14'b10110100001111: oled_data = 16'b1111111111111111;
				14'b10110110001111: oled_data = 16'b1111111111111111;
				14'b10111000001111: oled_data = 16'b1111111111111111;
				14'b10111010001111: oled_data = 16'b1111111111111111;
				14'b10111100001111: oled_data = 16'b1111111111111111;
				14'b10111110001111: oled_data = 16'b1111111111111111;
				14'b00000000010000: oled_data = 16'b1111111111111111;
				14'b00000010010000: oled_data = 16'b1111111111111111;
				14'b00000100010000: oled_data = 16'b1111111111111111;
				14'b00000110010000: oled_data = 16'b1111111111111111;
				14'b00001000010000: oled_data = 16'b1111111111111111;
				14'b00001010010000: oled_data = 16'b1111111111111111;
				14'b00001100010000: oled_data = 16'b1111111111111111;
				14'b00001110010000: oled_data = 16'b1111111111111111;
				14'b00010000010000: oled_data = 16'b1111111111111111;
				14'b00010010010000: oled_data = 16'b1111111111111111;
				14'b00010100010000: oled_data = 16'b1111111111111111;
				14'b00010110010000: oled_data = 16'b1111111111111111;
				14'b00011000010000: oled_data = 16'b1111111111111111;
				14'b00011010010000: oled_data = 16'b1111111111111111;
				14'b00011100010000: oled_data = 16'b1111111111111111;
				14'b00011110010000: oled_data = 16'b1111111111111111;
				14'b00100000010000: oled_data = 16'b1111111111111111;
				14'b00100010010000: oled_data = 16'b1111111111111111;
				14'b00100100010000: oled_data = 16'b1111111111111111;
				14'b00100110010000: oled_data = 16'b1111111111111111;
				14'b00101000010000: oled_data = 16'b1111011111011110;
				14'b00101010010000: oled_data = 16'b1000010010010011;
				14'b00101100010000: oled_data = 16'b1110011100111100;
				14'b00101110010000: oled_data = 16'b1111111111111111;
				14'b00110000010000: oled_data = 16'b1000110010110100;
				14'b00110010010000: oled_data = 16'b1010110110110111;
				14'b00110100010000: oled_data = 16'b1111111111111111;
				14'b00110110010000: oled_data = 16'b1101011011111011;
				14'b00111000010000: oled_data = 16'b1000110010110100;
				14'b00111010010000: oled_data = 16'b1110111101111101;
				14'b00111100010000: oled_data = 16'b0111110001010010;
				14'b00111110010000: oled_data = 16'b1111011110111110;
				14'b01000000010000: oled_data = 16'b1111111111111111;
				14'b01000010010000: oled_data = 16'b1111111111111111;
				14'b01000100010000: oled_data = 16'b1101111100111100;
				14'b01000110010000: oled_data = 16'b0111110001010010;
				14'b01001000010000: oled_data = 16'b1110111101111101;
				14'b01001010010000: oled_data = 16'b1000010001110011;
				14'b01001100010000: oled_data = 16'b1111011110111110;
				14'b01001110010000: oled_data = 16'b1101011011011011;
				14'b01010000010000: oled_data = 16'b1000110011010100;
				14'b01010010010000: oled_data = 16'b1111111111111111;
				14'b01010100010000: oled_data = 16'b1111111111111111;
				14'b01010110010000: oled_data = 16'b1101011011011011;
				14'b01011000010000: oled_data = 16'b0110001110110000;
				14'b01011010010000: oled_data = 16'b1110011101011101;
				14'b01011100010000: oled_data = 16'b1111111111111111;
				14'b01011110010000: oled_data = 16'b1111111111111111;
				14'b01100000010000: oled_data = 16'b1110111110011101;
				14'b01100010010000: oled_data = 16'b1000010001110011;
				14'b01100100010000: oled_data = 16'b1111011110111110;
				14'b01100110010000: oled_data = 16'b1111011111011110;
				14'b01101000010000: oled_data = 16'b0111010000110010;
				14'b01101010010000: oled_data = 16'b1100011001111010;
				14'b01101100010000: oled_data = 16'b1111111111111111;
				14'b01101110010000: oled_data = 16'b1100011001011001;
				14'b01110000010000: oled_data = 16'b1001110100110101;
				14'b01110010010000: oled_data = 16'b1111111111111111;
				14'b01110100010000: oled_data = 16'b1011010111111000;
				14'b01110110010000: oled_data = 16'b0110001110010000;
				14'b01111000010000: oled_data = 16'b0111010000010001;
				14'b01111010010000: oled_data = 16'b0110101111110001;
				14'b01111100010000: oled_data = 16'b1011111000011000;
				14'b01111110010000: oled_data = 16'b1111011110111110;
				14'b10000000010000: oled_data = 16'b1000010001110011;
				14'b10000010010000: oled_data = 16'b1110111110011110;
				14'b10000100010000: oled_data = 16'b1111111111111111;
				14'b10000110010000: oled_data = 16'b1110111110011101;
				14'b10001000010000: oled_data = 16'b0110101111010001;
				14'b10001010010000: oled_data = 16'b1100011001111010;
				14'b10001100010000: oled_data = 16'b1111111111111111;
				14'b10001110010000: oled_data = 16'b1110011101011100;
				14'b10010000010000: oled_data = 16'b0111110000110010;
				14'b10010010010000: oled_data = 16'b0111001111110001;
				14'b10010100010000: oled_data = 16'b0110101111110001;
				14'b10010110010000: oled_data = 16'b1010110110110111;
				14'b10011000010000: oled_data = 16'b1111111111111111;
				14'b10011010010000: oled_data = 16'b1111111111111111;
				14'b10011100010000: oled_data = 16'b1111111111111111;
				14'b10011110010000: oled_data = 16'b1111111111111111;
				14'b10100000010000: oled_data = 16'b1111011110111110;
				14'b10100010010000: oled_data = 16'b1110111110011101;
				14'b10100100010000: oled_data = 16'b1101011100111011;
				14'b10100110010000: oled_data = 16'b1100111011111010;
				14'b10101000010000: oled_data = 16'b1100111100011010;
				14'b10101010010000: oled_data = 16'b1101111101011011;
				14'b10101100010000: oled_data = 16'b1101111101011011;
				14'b10101110010000: oled_data = 16'b1101111101011011;
				14'b10110000010000: oled_data = 16'b1110011101111100;
				14'b10110010010000: oled_data = 16'b1110111110111101;
				14'b10110100010000: oled_data = 16'b1111111111111111;
				14'b10110110010000: oled_data = 16'b1111111111111111;
				14'b10111000010000: oled_data = 16'b1111111111111111;
				14'b10111010010000: oled_data = 16'b1111111111111111;
				14'b10111100010000: oled_data = 16'b1111111111111111;
				14'b10111110010000: oled_data = 16'b1111111111111111;
				14'b00000000010001: oled_data = 16'b1111111111111111;
				14'b00000010010001: oled_data = 16'b1111111111111111;
				14'b00000100010001: oled_data = 16'b1111111111111111;
				14'b00000110010001: oled_data = 16'b1111111111111111;
				14'b00001000010001: oled_data = 16'b1111111111111111;
				14'b00001010010001: oled_data = 16'b1111111111111111;
				14'b00001100010001: oled_data = 16'b1111111111111111;
				14'b00001110010001: oled_data = 16'b1111111111111111;
				14'b00010000010001: oled_data = 16'b1111111111111111;
				14'b00010010010001: oled_data = 16'b1111111111111111;
				14'b00010100010001: oled_data = 16'b1111111111111111;
				14'b00010110010001: oled_data = 16'b1111111111111111;
				14'b00011000010001: oled_data = 16'b1111111111111111;
				14'b00011010010001: oled_data = 16'b1111111111111111;
				14'b00011100010001: oled_data = 16'b1111111111111111;
				14'b00011110010001: oled_data = 16'b1111111111111111;
				14'b00100000010001: oled_data = 16'b1111111111111111;
				14'b00100010010001: oled_data = 16'b1111111111111111;
				14'b00100100010001: oled_data = 16'b1111111111111111;
				14'b00100110010001: oled_data = 16'b1111111111111111;
				14'b00101000010001: oled_data = 16'b1111111111111111;
				14'b00101010010001: oled_data = 16'b1111011111011110;
				14'b00101100010001: oled_data = 16'b1111011111011110;
				14'b00101110010001: oled_data = 16'b1111111111111111;
				14'b00110000010001: oled_data = 16'b1111011111011110;
				14'b00110010010001: oled_data = 16'b1111111111111111;
				14'b00110100010001: oled_data = 16'b1111111111111111;
				14'b00110110010001: oled_data = 16'b1111011111011110;
				14'b00111000010001: oled_data = 16'b1111011111011110;
				14'b00111010010001: oled_data = 16'b1111011111011110;
				14'b00111100010001: oled_data = 16'b1111011111011110;
				14'b00111110010001: oled_data = 16'b1111111111111111;
				14'b01000000010001: oled_data = 16'b1111111111111111;
				14'b01000010010001: oled_data = 16'b1111111111111111;
				14'b01000100010001: oled_data = 16'b1111111111111111;
				14'b01000110010001: oled_data = 16'b1111011110111110;
				14'b01001000010001: oled_data = 16'b1111011111011110;
				14'b01001010010001: oled_data = 16'b1111011111011110;
				14'b01001100010001: oled_data = 16'b1111111111111111;
				14'b01001110010001: oled_data = 16'b1111011111011110;
				14'b01010000010001: oled_data = 16'b1111011111011110;
				14'b01010010010001: oled_data = 16'b1111111111111111;
				14'b01010100010001: oled_data = 16'b1111111111111111;
				14'b01010110010001: oled_data = 16'b1111111111111111;
				14'b01011000010001: oled_data = 16'b1111011111011110;
				14'b01011010010001: oled_data = 16'b1111111111111111;
				14'b01011100010001: oled_data = 16'b1111111111111111;
				14'b01011110010001: oled_data = 16'b1111111111111111;
				14'b01100000010001: oled_data = 16'b1111111111111111;
				14'b01100010010001: oled_data = 16'b1111011111011110;
				14'b01100100010001: oled_data = 16'b1111111111111111;
				14'b01100110010001: oled_data = 16'b1111111111111111;
				14'b01101000010001: oled_data = 16'b1111011111011110;
				14'b01101010010001: oled_data = 16'b1111111111111111;
				14'b01101100010001: oled_data = 16'b1111111111111111;
				14'b01101110010001: oled_data = 16'b1111011111011110;
				14'b01110000010001: oled_data = 16'b1111011111011110;
				14'b01110010010001: oled_data = 16'b1111111111111111;
				14'b01110100010001: oled_data = 16'b1111011111011110;
				14'b01110110010001: oled_data = 16'b1111011110111110;
				14'b01111000010001: oled_data = 16'b1110111110011110;
				14'b01111010010001: oled_data = 16'b1110111110011110;
				14'b01111100010001: oled_data = 16'b1111011111011110;
				14'b01111110010001: oled_data = 16'b1111111111111111;
				14'b10000000010001: oled_data = 16'b1111011111011110;
				14'b10000010010001: oled_data = 16'b1111111111111111;
				14'b10000100010001: oled_data = 16'b1111111111111111;
				14'b10000110010001: oled_data = 16'b1111111111111111;
				14'b10001000010001: oled_data = 16'b1111011111011110;
				14'b10001010010001: oled_data = 16'b1111011111011110;
				14'b10001100010001: oled_data = 16'b1111111111111111;
				14'b10001110010001: oled_data = 16'b1111111111111111;
				14'b10010000010001: oled_data = 16'b1111111111111111;
				14'b10010010010001: oled_data = 16'b1110011101111101;
				14'b10010100010001: oled_data = 16'b1111011110111110;
				14'b10010110010001: oled_data = 16'b1111111111111111;
				14'b10011000010001: oled_data = 16'b1111111111111111;
				14'b10011010010001: oled_data = 16'b1111111111111111;
				14'b10011100010001: oled_data = 16'b1111111111111111;
				14'b10011110010001: oled_data = 16'b1111111111111111;
				14'b10100000010001: oled_data = 16'b1111011111111111;
				14'b10100010010001: oled_data = 16'b1110111110111101;
				14'b10100100010001: oled_data = 16'b1110011101111100;
				14'b10100110010001: oled_data = 16'b1100111100011010;
				14'b10101000010001: oled_data = 16'b1100111100011010;
				14'b10101010010001: oled_data = 16'b1101011100111010;
				14'b10101100010001: oled_data = 16'b1101111101011011;
				14'b10101110010001: oled_data = 16'b1101111101011011;
				14'b10110000010001: oled_data = 16'b1101111101011011;
				14'b10110010010001: oled_data = 16'b1110011101111100;
				14'b10110100010001: oled_data = 16'b1110111110111110;
				14'b10110110010001: oled_data = 16'b1111111111111111;
				14'b10111000010001: oled_data = 16'b1111111111111111;
				14'b10111010010001: oled_data = 16'b1111111111111111;
				14'b10111100010001: oled_data = 16'b1111111111111111;
				14'b10111110010001: oled_data = 16'b1111111111111111;
				14'b00000000010010: oled_data = 16'b1111111111111111;
				14'b00000010010010: oled_data = 16'b1111111111111111;
				14'b00000100010010: oled_data = 16'b1111111111111111;
				14'b00000110010010: oled_data = 16'b1111111111111111;
				14'b00001000010010: oled_data = 16'b1111111111111111;
				14'b00001010010010: oled_data = 16'b1111111111111111;
				14'b00001100010010: oled_data = 16'b1111111111111111;
				14'b00001110010010: oled_data = 16'b1111111111111111;
				14'b00010000010010: oled_data = 16'b1111111111111111;
				14'b00010010010010: oled_data = 16'b1111111111111111;
				14'b00010100010010: oled_data = 16'b1111111111111111;
				14'b00010110010010: oled_data = 16'b1111111111111111;
				14'b00011000010010: oled_data = 16'b1111111111111111;
				14'b00011010010010: oled_data = 16'b1111111111111111;
				14'b00011100010010: oled_data = 16'b1111111111111111;
				14'b00011110010010: oled_data = 16'b1111111111111111;
				14'b00100000010010: oled_data = 16'b1111111111111111;
				14'b00100010010010: oled_data = 16'b1111111111111111;
				14'b00100100010010: oled_data = 16'b1111111111111111;
				14'b00100110010010: oled_data = 16'b1111111111111111;
				14'b00101000010010: oled_data = 16'b1111111111111111;
				14'b00101010010010: oled_data = 16'b1111111111111111;
				14'b00101100010010: oled_data = 16'b1111111111111111;
				14'b00101110010010: oled_data = 16'b1111111111111111;
				14'b00110000010010: oled_data = 16'b1111111111111111;
				14'b00110010010010: oled_data = 16'b1111111111111111;
				14'b00110100010010: oled_data = 16'b1111111111111111;
				14'b00110110010010: oled_data = 16'b1111111111111111;
				14'b00111000010010: oled_data = 16'b1111111111111111;
				14'b00111010010010: oled_data = 16'b1111111111111111;
				14'b00111100010010: oled_data = 16'b1111111111111111;
				14'b00111110010010: oled_data = 16'b1111111111111111;
				14'b01000000010010: oled_data = 16'b1111111111111111;
				14'b01000010010010: oled_data = 16'b1111111111111111;
				14'b01000100010010: oled_data = 16'b1111111111111111;
				14'b01000110010010: oled_data = 16'b1111111111111111;
				14'b01001000010010: oled_data = 16'b1111111111111111;
				14'b01001010010010: oled_data = 16'b1111111111111111;
				14'b01001100010010: oled_data = 16'b1111111111111111;
				14'b01001110010010: oled_data = 16'b1111111111111111;
				14'b01010000010010: oled_data = 16'b1111111111111111;
				14'b01010010010010: oled_data = 16'b1111111111111111;
				14'b01010100010010: oled_data = 16'b1111111111111111;
				14'b01010110010010: oled_data = 16'b1111111111111111;
				14'b01011000010010: oled_data = 16'b1111111111111111;
				14'b01011010010010: oled_data = 16'b1111111111111111;
				14'b01011100010010: oled_data = 16'b1111111111111111;
				14'b01011110010010: oled_data = 16'b1111111111111111;
				14'b01100000010010: oled_data = 16'b1111111111111111;
				14'b01100010010010: oled_data = 16'b1111111111111111;
				14'b01100100010010: oled_data = 16'b1111111111111111;
				14'b01100110010010: oled_data = 16'b1111111111111111;
				14'b01101000010010: oled_data = 16'b1111111111111111;
				14'b01101010010010: oled_data = 16'b1111111111111111;
				14'b01101100010010: oled_data = 16'b1111111111111111;
				14'b01101110010010: oled_data = 16'b1111111111111111;
				14'b01110000010010: oled_data = 16'b1111111111111111;
				14'b01110010010010: oled_data = 16'b1111111111111111;
				14'b01110100010010: oled_data = 16'b1111111111111111;
				14'b01110110010010: oled_data = 16'b1111111111111111;
				14'b01111000010010: oled_data = 16'b1111111111111111;
				14'b01111010010010: oled_data = 16'b1111111111111111;
				14'b01111100010010: oled_data = 16'b1111111111111111;
				14'b01111110010010: oled_data = 16'b1111111111111111;
				14'b10000000010010: oled_data = 16'b1111111111111111;
				14'b10000010010010: oled_data = 16'b1111111111111111;
				14'b10000100010010: oled_data = 16'b1111111111111111;
				14'b10000110010010: oled_data = 16'b1111111111111111;
				14'b10001000010010: oled_data = 16'b1111111111111111;
				14'b10001010010010: oled_data = 16'b1111111111111111;
				14'b10001100010010: oled_data = 16'b1111111111111111;
				14'b10001110010010: oled_data = 16'b1111111111111111;
				14'b10010000010010: oled_data = 16'b1111111111111111;
				14'b10010010010010: oled_data = 16'b1111111111111111;
				14'b10010100010010: oled_data = 16'b1111111111111111;
				14'b10010110010010: oled_data = 16'b1111111111111111;
				14'b10011000010010: oled_data = 16'b1111111111111111;
				14'b10011010010010: oled_data = 16'b1111111111111111;
				14'b10011100010010: oled_data = 16'b1111111111111111;
				14'b10011110010010: oled_data = 16'b1111111111111111;
				14'b10100000010010: oled_data = 16'b1111111111111111;
				14'b10100010010010: oled_data = 16'b1111011111011110;
				14'b10100100010010: oled_data = 16'b1110111110111101;
				14'b10100110010010: oled_data = 16'b1101111101011011;
				14'b10101000010010: oled_data = 16'b1100111011111001;
				14'b10101010010010: oled_data = 16'b1101011100011010;
				14'b10101100010010: oled_data = 16'b1101011100111011;
				14'b10101110010010: oled_data = 16'b1101111101011011;
				14'b10110000010010: oled_data = 16'b1101111101011011;
				14'b10110010010010: oled_data = 16'b1101111101011011;
				14'b10110100010010: oled_data = 16'b1110011101111100;
				14'b10110110010010: oled_data = 16'b1110111110111110;
				14'b10111000010010: oled_data = 16'b1111011111111110;
				14'b10111010010010: oled_data = 16'b1111111111111111;
				14'b10111100010010: oled_data = 16'b1111111111111111;
				14'b10111110010010: oled_data = 16'b1111111111111111;
				14'b00000000010011: oled_data = 16'b1111111111111111;
				14'b00000010010011: oled_data = 16'b1111111111111111;
				14'b00000100010011: oled_data = 16'b1111111111111111;
				14'b00000110010011: oled_data = 16'b1111111111111111;
				14'b00001000010011: oled_data = 16'b1111111111111111;
				14'b00001010010011: oled_data = 16'b1111111111111111;
				14'b00001100010011: oled_data = 16'b1111111111111111;
				14'b00001110010011: oled_data = 16'b1111111111111111;
				14'b00010000010011: oled_data = 16'b1111111111111111;
				14'b00010010010011: oled_data = 16'b1111111111111111;
				14'b00010100010011: oled_data = 16'b1111111111111111;
				14'b00010110010011: oled_data = 16'b1111111111111111;
				14'b00011000010011: oled_data = 16'b1111111111111111;
				14'b00011010010011: oled_data = 16'b1111111111111111;
				14'b00011100010011: oled_data = 16'b1111111111111111;
				14'b00011110010011: oled_data = 16'b1111111111111111;
				14'b00100000010011: oled_data = 16'b1111111111111111;
				14'b00100010010011: oled_data = 16'b1111111111111111;
				14'b00100100010011: oled_data = 16'b1111111111111111;
				14'b00100110010011: oled_data = 16'b1111111111111111;
				14'b00101000010011: oled_data = 16'b1111111111111111;
				14'b00101010010011: oled_data = 16'b1111111111111111;
				14'b00101100010011: oled_data = 16'b1111111111111111;
				14'b00101110010011: oled_data = 16'b1111111111111111;
				14'b00110000010011: oled_data = 16'b1111111111111111;
				14'b00110010010011: oled_data = 16'b1111111111111111;
				14'b00110100010011: oled_data = 16'b1111111111111111;
				14'b00110110010011: oled_data = 16'b1111111111111111;
				14'b00111000010011: oled_data = 16'b1111111111111111;
				14'b00111010010011: oled_data = 16'b1111111111111111;
				14'b00111100010011: oled_data = 16'b1111111111111111;
				14'b00111110010011: oled_data = 16'b1111111111111111;
				14'b01000000010011: oled_data = 16'b1111111111111111;
				14'b01000010010011: oled_data = 16'b1111111111111111;
				14'b01000100010011: oled_data = 16'b1111111111111111;
				14'b01000110010011: oled_data = 16'b1111111111111111;
				14'b01001000010011: oled_data = 16'b1111111111111111;
				14'b01001010010011: oled_data = 16'b1111111111111111;
				14'b01001100010011: oled_data = 16'b1111111111111111;
				14'b01001110010011: oled_data = 16'b1111111111111111;
				14'b01010000010011: oled_data = 16'b1111111111111111;
				14'b01010010010011: oled_data = 16'b1111111111111111;
				14'b01010100010011: oled_data = 16'b1111111111111111;
				14'b01010110010011: oled_data = 16'b1111111111111111;
				14'b01011000010011: oled_data = 16'b1111111111111111;
				14'b01011010010011: oled_data = 16'b1111111111111111;
				14'b01011100010011: oled_data = 16'b1111111111111111;
				14'b01011110010011: oled_data = 16'b1111111111111111;
				14'b01100000010011: oled_data = 16'b1111111111111111;
				14'b01100010010011: oled_data = 16'b1111111111111111;
				14'b01100100010011: oled_data = 16'b1111111111111111;
				14'b01100110010011: oled_data = 16'b1111111111111111;
				14'b01101000010011: oled_data = 16'b1111111111111111;
				14'b01101010010011: oled_data = 16'b1111111111111111;
				14'b01101100010011: oled_data = 16'b1111111111111111;
				14'b01101110010011: oled_data = 16'b1111111111111111;
				14'b01110000010011: oled_data = 16'b1111111111111111;
				14'b01110010010011: oled_data = 16'b1111111111111111;
				14'b01110100010011: oled_data = 16'b1111111111111111;
				14'b01110110010011: oled_data = 16'b1111111111111111;
				14'b01111000010011: oled_data = 16'b1111111111111111;
				14'b01111010010011: oled_data = 16'b1111111111111111;
				14'b01111100010011: oled_data = 16'b1111111111111111;
				14'b01111110010011: oled_data = 16'b1111111111111111;
				14'b10000000010011: oled_data = 16'b1111111111111111;
				14'b10000010010011: oled_data = 16'b1111111111111111;
				14'b10000100010011: oled_data = 16'b1111111111111111;
				14'b10000110010011: oled_data = 16'b1111111111111111;
				14'b10001000010011: oled_data = 16'b1111111111111111;
				14'b10001010010011: oled_data = 16'b1111111111111111;
				14'b10001100010011: oled_data = 16'b1111111111111111;
				14'b10001110010011: oled_data = 16'b1111111111111111;
				14'b10010000010011: oled_data = 16'b1111111111111111;
				14'b10010010010011: oled_data = 16'b1111111111111111;
				14'b10010100010011: oled_data = 16'b1111111111111111;
				14'b10010110010011: oled_data = 16'b1111111111111111;
				14'b10011000010011: oled_data = 16'b1111111111111111;
				14'b10011010010011: oled_data = 16'b1111111111111111;
				14'b10011100010011: oled_data = 16'b1111111111111111;
				14'b10011110010011: oled_data = 16'b1111111111111111;
				14'b10100000010011: oled_data = 16'b1111111111111111;
				14'b10100010010011: oled_data = 16'b1111111111111111;
				14'b10100100010011: oled_data = 16'b1111011111011110;
				14'b10100110010011: oled_data = 16'b1110111110011101;
				14'b10101000010011: oled_data = 16'b1101011101011010;
				14'b10101010010011: oled_data = 16'b1100111100011001;
				14'b10101100010011: oled_data = 16'b1101011100011010;
				14'b10101110010011: oled_data = 16'b1101111101011011;
				14'b10110000010011: oled_data = 16'b1101111101011011;
				14'b10110010010011: oled_data = 16'b1101111101011011;
				14'b10110100010011: oled_data = 16'b1101111101011011;
				14'b10110110010011: oled_data = 16'b1110011101111100;
				14'b10111000010011: oled_data = 16'b1110111110111101;
				14'b10111010010011: oled_data = 16'b1111011111011110;
				14'b10111100010011: oled_data = 16'b1111111111111111;
				14'b10111110010011: oled_data = 16'b1111111111111111;
				14'b00000000010100: oled_data = 16'b1111111111111111;
				14'b00000010010100: oled_data = 16'b1111111111111111;
				14'b00000100010100: oled_data = 16'b1111111111111111;
				14'b00000110010100: oled_data = 16'b1111111111111111;
				14'b00001000010100: oled_data = 16'b1111111111111111;
				14'b00001010010100: oled_data = 16'b1111111111111111;
				14'b00001100010100: oled_data = 16'b1111111111111111;
				14'b00001110010100: oled_data = 16'b1111111111111111;
				14'b00010000010100: oled_data = 16'b1111111111111111;
				14'b00010010010100: oled_data = 16'b1111111111111111;
				14'b00010100010100: oled_data = 16'b1111111111111111;
				14'b00010110010100: oled_data = 16'b1111111111111111;
				14'b00011000010100: oled_data = 16'b1111111111111111;
				14'b00011010010100: oled_data = 16'b1111111111111111;
				14'b00011100010100: oled_data = 16'b1111111111111111;
				14'b00011110010100: oled_data = 16'b1111111111111111;
				14'b00100000010100: oled_data = 16'b1111111111111111;
				14'b00100010010100: oled_data = 16'b1111111111111111;
				14'b00100100010100: oled_data = 16'b1111111111111111;
				14'b00100110010100: oled_data = 16'b1111111111111111;
				14'b00101000010100: oled_data = 16'b1111111111111111;
				14'b00101010010100: oled_data = 16'b1111111111111111;
				14'b00101100010100: oled_data = 16'b1111111111111111;
				14'b00101110010100: oled_data = 16'b1111111111111111;
				14'b00110000010100: oled_data = 16'b1111111111111111;
				14'b00110010010100: oled_data = 16'b1111111111111111;
				14'b00110100010100: oled_data = 16'b1111111111111111;
				14'b00110110010100: oled_data = 16'b1111111111111111;
				14'b00111000010100: oled_data = 16'b1111111111111111;
				14'b00111010010100: oled_data = 16'b1111111111111111;
				14'b00111100010100: oled_data = 16'b1111111111111111;
				14'b00111110010100: oled_data = 16'b1111111111111111;
				14'b01000000010100: oled_data = 16'b1111111111111111;
				14'b01000010010100: oled_data = 16'b1111111111111111;
				14'b01000100010100: oled_data = 16'b1111111111111111;
				14'b01000110010100: oled_data = 16'b1111111111111111;
				14'b01001000010100: oled_data = 16'b1111111111111111;
				14'b01001010010100: oled_data = 16'b1111111111111111;
				14'b01001100010100: oled_data = 16'b1111111111111111;
				14'b01001110010100: oled_data = 16'b1111111111111111;
				14'b01010000010100: oled_data = 16'b1111111111111111;
				14'b01010010010100: oled_data = 16'b1111111111111111;
				14'b01010100010100: oled_data = 16'b1111111111111111;
				14'b01010110010100: oled_data = 16'b1111111111111111;
				14'b01011000010100: oled_data = 16'b1111111111111111;
				14'b01011010010100: oled_data = 16'b1111111111111111;
				14'b01011100010100: oled_data = 16'b1111111111111111;
				14'b01011110010100: oled_data = 16'b1111111111111111;
				14'b01100000010100: oled_data = 16'b1111111111111111;
				14'b01100010010100: oled_data = 16'b1111111111111111;
				14'b01100100010100: oled_data = 16'b1111111111111111;
				14'b01100110010100: oled_data = 16'b1111111111111111;
				14'b01101000010100: oled_data = 16'b1111111111111111;
				14'b01101010010100: oled_data = 16'b1111111111111111;
				14'b01101100010100: oled_data = 16'b1111111111111111;
				14'b01101110010100: oled_data = 16'b1111111111111111;
				14'b01110000010100: oled_data = 16'b1111111111111111;
				14'b01110010010100: oled_data = 16'b1111111111111111;
				14'b01110100010100: oled_data = 16'b1111111111111111;
				14'b01110110010100: oled_data = 16'b1111111111111111;
				14'b01111000010100: oled_data = 16'b1111111111111111;
				14'b01111010010100: oled_data = 16'b1111111111111111;
				14'b01111100010100: oled_data = 16'b1111111111111111;
				14'b01111110010100: oled_data = 16'b1111111111111111;
				14'b10000000010100: oled_data = 16'b1111111111111111;
				14'b10000010010100: oled_data = 16'b1111111111111111;
				14'b10000100010100: oled_data = 16'b1111111111111111;
				14'b10000110010100: oled_data = 16'b1111111111111111;
				14'b10001000010100: oled_data = 16'b1111111111111111;
				14'b10001010010100: oled_data = 16'b1111111111111111;
				14'b10001100010100: oled_data = 16'b1111111111111111;
				14'b10001110010100: oled_data = 16'b1111111111111111;
				14'b10010000010100: oled_data = 16'b1111111111111111;
				14'b10010010010100: oled_data = 16'b1111111111111111;
				14'b10010100010100: oled_data = 16'b1111111111111111;
				14'b10010110010100: oled_data = 16'b1111111111111111;
				14'b10011000010100: oled_data = 16'b1111111111111111;
				14'b10011010010100: oled_data = 16'b1111111111111111;
				14'b10011100010100: oled_data = 16'b1111111111111111;
				14'b10011110010100: oled_data = 16'b1111111111111111;
				14'b10100000010100: oled_data = 16'b1111111111111111;
				14'b10100010010100: oled_data = 16'b1111111111111111;
				14'b10100100010100: oled_data = 16'b1111111111111111;
				14'b10100110010100: oled_data = 16'b1111011111011110;
				14'b10101000010100: oled_data = 16'b1110011110011100;
				14'b10101010010100: oled_data = 16'b1101011100111010;
				14'b10101100010100: oled_data = 16'b1100111100011001;
				14'b10101110010100: oled_data = 16'b1101011100111010;
				14'b10110000010100: oled_data = 16'b1101111101011011;
				14'b10110010010100: oled_data = 16'b1101111101011011;
				14'b10110100010100: oled_data = 16'b1101111101011011;
				14'b10110110010100: oled_data = 16'b1101111101011011;
				14'b10111000010100: oled_data = 16'b1110011101111100;
				14'b10111010010100: oled_data = 16'b1110111110011101;
				14'b10111100010100: oled_data = 16'b1111011111011110;
				14'b10111110010100: oled_data = 16'b1111111111111111;
				14'b00000000010101: oled_data = 16'b1111111111111111;
				14'b00000010010101: oled_data = 16'b1111111111111111;
				14'b00000100010101: oled_data = 16'b1111111111111111;
				14'b00000110010101: oled_data = 16'b1111111111111111;
				14'b00001000010101: oled_data = 16'b1111111111111111;
				14'b00001010010101: oled_data = 16'b1111111111111111;
				14'b00001100010101: oled_data = 16'b1111111111111111;
				14'b00001110010101: oled_data = 16'b1111111111111111;
				14'b00010000010101: oled_data = 16'b1111111111111111;
				14'b00010010010101: oled_data = 16'b1111111111111111;
				14'b00010100010101: oled_data = 16'b1111111111111111;
				14'b00010110010101: oled_data = 16'b1111111111111111;
				14'b00011000010101: oled_data = 16'b1111111111111111;
				14'b00011010010101: oled_data = 16'b1111111111111111;
				14'b00011100010101: oled_data = 16'b1111111111111111;
				14'b00011110010101: oled_data = 16'b1111111111111111;
				14'b00100000010101: oled_data = 16'b1111111111111111;
				14'b00100010010101: oled_data = 16'b1111111111111111;
				14'b00100100010101: oled_data = 16'b1111111111111111;
				14'b00100110010101: oled_data = 16'b1111111111111111;
				14'b00101000010101: oled_data = 16'b1111111111111111;
				14'b00101010010101: oled_data = 16'b1111111111111111;
				14'b00101100010101: oled_data = 16'b1111111111111111;
				14'b00101110010101: oled_data = 16'b1111111111111111;
				14'b00110000010101: oled_data = 16'b1111111111111111;
				14'b00110010010101: oled_data = 16'b1111111111111111;
				14'b00110100010101: oled_data = 16'b1111111111111111;
				14'b00110110010101: oled_data = 16'b1111111111111111;
				14'b00111000010101: oled_data = 16'b1111111111111111;
				14'b00111010010101: oled_data = 16'b1111111111111111;
				14'b00111100010101: oled_data = 16'b1111111111111111;
				14'b00111110010101: oled_data = 16'b1111111111111111;
				14'b01000000010101: oled_data = 16'b1111111111111111;
				14'b01000010010101: oled_data = 16'b1111111111111111;
				14'b01000100010101: oled_data = 16'b1111111111111111;
				14'b01000110010101: oled_data = 16'b1111111111111111;
				14'b01001000010101: oled_data = 16'b1111111111111111;
				14'b01001010010101: oled_data = 16'b1111111111111111;
				14'b01001100010101: oled_data = 16'b1111111111111111;
				14'b01001110010101: oled_data = 16'b1111111111111111;
				14'b01010000010101: oled_data = 16'b1111111111111111;
				14'b01010010010101: oled_data = 16'b1111111111111111;
				14'b01010100010101: oled_data = 16'b1111111111111111;
				14'b01010110010101: oled_data = 16'b1111111111111111;
				14'b01011000010101: oled_data = 16'b1111111111111111;
				14'b01011010010101: oled_data = 16'b1111111111111111;
				14'b01011100010101: oled_data = 16'b1111111111111111;
				14'b01011110010101: oled_data = 16'b1111111111111111;
				14'b01100000010101: oled_data = 16'b1111111111111111;
				14'b01100010010101: oled_data = 16'b1111111111111111;
				14'b01100100010101: oled_data = 16'b1111111111111111;
				14'b01100110010101: oled_data = 16'b1111111111111111;
				14'b01101000010101: oled_data = 16'b1111111111111111;
				14'b01101010010101: oled_data = 16'b1111111111111111;
				14'b01101100010101: oled_data = 16'b1111111111111111;
				14'b01101110010101: oled_data = 16'b1111111111111111;
				14'b01110000010101: oled_data = 16'b1111111111111111;
				14'b01110010010101: oled_data = 16'b1111111111111111;
				14'b01110100010101: oled_data = 16'b1111111111111111;
				14'b01110110010101: oled_data = 16'b1111111111111111;
				14'b01111000010101: oled_data = 16'b1111111111111111;
				14'b01111010010101: oled_data = 16'b1111111111111111;
				14'b01111100010101: oled_data = 16'b1111111111111111;
				14'b01111110010101: oled_data = 16'b1111111111111111;
				14'b10000000010101: oled_data = 16'b1111111111111111;
				14'b10000010010101: oled_data = 16'b1111111111111111;
				14'b10000100010101: oled_data = 16'b1111111111111111;
				14'b10000110010101: oled_data = 16'b1111111111111111;
				14'b10001000010101: oled_data = 16'b1111111111111111;
				14'b10001010010101: oled_data = 16'b1111111111111111;
				14'b10001100010101: oled_data = 16'b1111111111111111;
				14'b10001110010101: oled_data = 16'b1111111111111111;
				14'b10010000010101: oled_data = 16'b1111111111111111;
				14'b10010010010101: oled_data = 16'b1111111111111111;
				14'b10010100010101: oled_data = 16'b1111111111111111;
				14'b10010110010101: oled_data = 16'b1111111111111111;
				14'b10011000010101: oled_data = 16'b1111111111111111;
				14'b10011010010101: oled_data = 16'b1111111111111111;
				14'b10011100010101: oled_data = 16'b1111111111111111;
				14'b10011110010101: oled_data = 16'b1111111111111111;
				14'b10100000010101: oled_data = 16'b1111111111111111;
				14'b10100010010101: oled_data = 16'b1111111111111111;
				14'b10100100010101: oled_data = 16'b1111111111111111;
				14'b10100110010101: oled_data = 16'b1111111111111111;
				14'b10101000010101: oled_data = 16'b1111011111011110;
				14'b10101010010101: oled_data = 16'b1110011110011100;
				14'b10101100010101: oled_data = 16'b1100111100011001;
				14'b10101110010101: oled_data = 16'b1100111100011001;
				14'b10110000010101: oled_data = 16'b1101011100111010;
				14'b10110010010101: oled_data = 16'b1101111101011011;
				14'b10110100010101: oled_data = 16'b1101111101011011;
				14'b10110110010101: oled_data = 16'b1101111101011011;
				14'b10111000010101: oled_data = 16'b1101111101011011;
				14'b10111010010101: oled_data = 16'b1101111101011011;
				14'b10111100010101: oled_data = 16'b1110011110011100;
				14'b10111110010101: oled_data = 16'b1110111110111101;
				14'b00000000010110: oled_data = 16'b1111111111111111;
				14'b00000010010110: oled_data = 16'b1111111111111111;
				14'b00000100010110: oled_data = 16'b1111111111111111;
				14'b00000110010110: oled_data = 16'b1111111111111111;
				14'b00001000010110: oled_data = 16'b1111111111111111;
				14'b00001010010110: oled_data = 16'b1111111111111111;
				14'b00001100010110: oled_data = 16'b1111111111111111;
				14'b00001110010110: oled_data = 16'b1111111111111111;
				14'b00010000010110: oled_data = 16'b1111111111111111;
				14'b00010010010110: oled_data = 16'b1111111111111111;
				14'b00010100010110: oled_data = 16'b1111111111111111;
				14'b00010110010110: oled_data = 16'b1111111111111111;
				14'b00011000010110: oled_data = 16'b1111111111111111;
				14'b00011010010110: oled_data = 16'b1111111111111111;
				14'b00011100010110: oled_data = 16'b1111111111111111;
				14'b00011110010110: oled_data = 16'b1111111111111111;
				14'b00100000010110: oled_data = 16'b1111111111111111;
				14'b00100010010110: oled_data = 16'b1111111111111111;
				14'b00100100010110: oled_data = 16'b1111111111111111;
				14'b00100110010110: oled_data = 16'b1111111111111111;
				14'b00101000010110: oled_data = 16'b1111111111111111;
				14'b00101010010110: oled_data = 16'b1111111111111111;
				14'b00101100010110: oled_data = 16'b1111111111111111;
				14'b00101110010110: oled_data = 16'b1111111111111111;
				14'b00110000010110: oled_data = 16'b1111111111111111;
				14'b00110010010110: oled_data = 16'b1111111111111111;
				14'b00110100010110: oled_data = 16'b1111111111111111;
				14'b00110110010110: oled_data = 16'b1111111111111111;
				14'b00111000010110: oled_data = 16'b1111111111111111;
				14'b00111010010110: oled_data = 16'b1111111111111111;
				14'b00111100010110: oled_data = 16'b1111111111111111;
				14'b00111110010110: oled_data = 16'b1111111111111111;
				14'b01000000010110: oled_data = 16'b1111111111111111;
				14'b01000010010110: oled_data = 16'b1111111111111111;
				14'b01000100010110: oled_data = 16'b1111111111111111;
				14'b01000110010110: oled_data = 16'b1111111111111111;
				14'b01001000010110: oled_data = 16'b1111111111111111;
				14'b01001010010110: oled_data = 16'b1111111111111111;
				14'b01001100010110: oled_data = 16'b1111111111111111;
				14'b01001110010110: oled_data = 16'b1111111111111111;
				14'b01010000010110: oled_data = 16'b1111111111111111;
				14'b01010010010110: oled_data = 16'b1111111111111111;
				14'b01010100010110: oled_data = 16'b1111111111111111;
				14'b01010110010110: oled_data = 16'b1111111111111111;
				14'b01011000010110: oled_data = 16'b1111111111111111;
				14'b01011010010110: oled_data = 16'b1111111111111111;
				14'b01011100010110: oled_data = 16'b1111111111111111;
				14'b01011110010110: oled_data = 16'b1111111111111111;
				14'b01100000010110: oled_data = 16'b1111111111111111;
				14'b01100010010110: oled_data = 16'b1111111111111111;
				14'b01100100010110: oled_data = 16'b1111111111111111;
				14'b01100110010110: oled_data = 16'b1111111111111111;
				14'b01101000010110: oled_data = 16'b1111111111111111;
				14'b01101010010110: oled_data = 16'b1111111111111111;
				14'b01101100010110: oled_data = 16'b1111111111111111;
				14'b01101110010110: oled_data = 16'b1111111111111111;
				14'b01110000010110: oled_data = 16'b1111111111111111;
				14'b01110010010110: oled_data = 16'b1111111111111111;
				14'b01110100010110: oled_data = 16'b1111111111111111;
				14'b01110110010110: oled_data = 16'b1111111111111111;
				14'b01111000010110: oled_data = 16'b1111111111111111;
				14'b01111010010110: oled_data = 16'b1111111111111111;
				14'b01111100010110: oled_data = 16'b1111111111111111;
				14'b01111110010110: oled_data = 16'b1111111111111111;
				14'b10000000010110: oled_data = 16'b1111111111111111;
				14'b10000010010110: oled_data = 16'b1111111111111111;
				14'b10000100010110: oled_data = 16'b1111111111111111;
				14'b10000110010110: oled_data = 16'b1111111111111111;
				14'b10001000010110: oled_data = 16'b1111111111111111;
				14'b10001010010110: oled_data = 16'b1111111111111111;
				14'b10001100010110: oled_data = 16'b1111111111111111;
				14'b10001110010110: oled_data = 16'b1111111111111111;
				14'b10010000010110: oled_data = 16'b1111111111111111;
				14'b10010010010110: oled_data = 16'b1111111111111111;
				14'b10010100010110: oled_data = 16'b1111111111111111;
				14'b10010110010110: oled_data = 16'b1111111111111111;
				14'b10011000010110: oled_data = 16'b1111111111111111;
				14'b10011010010110: oled_data = 16'b1111111111111111;
				14'b10011100010110: oled_data = 16'b1111111111111111;
				14'b10011110010110: oled_data = 16'b1111111111111111;
				14'b10100000010110: oled_data = 16'b1111111111111111;
				14'b10100010010110: oled_data = 16'b1111111111111111;
				14'b10100100010110: oled_data = 16'b1111111111111111;
				14'b10100110010110: oled_data = 16'b1111111111111111;
				14'b10101000010110: oled_data = 16'b1111111111111111;
				14'b10101010010110: oled_data = 16'b1111011111011110;
				14'b10101100010110: oled_data = 16'b1110011101111100;
				14'b10101110010110: oled_data = 16'b1100111100011001;
				14'b10110000010110: oled_data = 16'b1100111100011001;
				14'b10110010010110: oled_data = 16'b1101011100111010;
				14'b10110100010110: oled_data = 16'b1101111101011011;
				14'b10110110010110: oled_data = 16'b1101111101011011;
				14'b10111000010110: oled_data = 16'b1101111101011011;
				14'b10111010010110: oled_data = 16'b1101111101011011;
				14'b10111100010110: oled_data = 16'b1101111101011011;
				14'b10111110010110: oled_data = 16'b1101111101111100;
				14'b00000000010111: oled_data = 16'b1111111111111111;
				14'b00000010010111: oled_data = 16'b1111111111111111;
				14'b00000100010111: oled_data = 16'b1111111111111111;
				14'b00000110010111: oled_data = 16'b1111111111111111;
				14'b00001000010111: oled_data = 16'b1111111111111111;
				14'b00001010010111: oled_data = 16'b1111111111111111;
				14'b00001100010111: oled_data = 16'b1111111111111111;
				14'b00001110010111: oled_data = 16'b1111111111111111;
				14'b00010000010111: oled_data = 16'b1111111111111111;
				14'b00010010010111: oled_data = 16'b1111111111111111;
				14'b00010100010111: oled_data = 16'b1111111111111111;
				14'b00010110010111: oled_data = 16'b1111111111111111;
				14'b00011000010111: oled_data = 16'b1111111111111111;
				14'b00011010010111: oled_data = 16'b1111111111111111;
				14'b00011100010111: oled_data = 16'b1111111111111111;
				14'b00011110010111: oled_data = 16'b1111111111111111;
				14'b00100000010111: oled_data = 16'b1111111111111111;
				14'b00100010010111: oled_data = 16'b1111111111111111;
				14'b00100100010111: oled_data = 16'b1111111111111111;
				14'b00100110010111: oled_data = 16'b1111111111111111;
				14'b00101000010111: oled_data = 16'b1111111111111111;
				14'b00101010010111: oled_data = 16'b1111111111111111;
				14'b00101100010111: oled_data = 16'b1111111111111111;
				14'b00101110010111: oled_data = 16'b1111111111111111;
				14'b00110000010111: oled_data = 16'b1111111111111111;
				14'b00110010010111: oled_data = 16'b1111111111111111;
				14'b00110100010111: oled_data = 16'b1111111111111111;
				14'b00110110010111: oled_data = 16'b1111111111111111;
				14'b00111000010111: oled_data = 16'b1111111111111111;
				14'b00111010010111: oled_data = 16'b1111111111111111;
				14'b00111100010111: oled_data = 16'b1111111111111111;
				14'b00111110010111: oled_data = 16'b1111111111111111;
				14'b01000000010111: oled_data = 16'b1111111111111111;
				14'b01000010010111: oled_data = 16'b1111111111111111;
				14'b01000100010111: oled_data = 16'b1111111111111111;
				14'b01000110010111: oled_data = 16'b1111111111111111;
				14'b01001000010111: oled_data = 16'b1111111111111111;
				14'b01001010010111: oled_data = 16'b1111111111111111;
				14'b01001100010111: oled_data = 16'b1111111111111111;
				14'b01001110010111: oled_data = 16'b1111111111111111;
				14'b01010000010111: oled_data = 16'b1111111111111111;
				14'b01010010010111: oled_data = 16'b1111111111111111;
				14'b01010100010111: oled_data = 16'b1111111111111111;
				14'b01010110010111: oled_data = 16'b1111111111111111;
				14'b01011000010111: oled_data = 16'b1111111111111111;
				14'b01011010010111: oled_data = 16'b1111111111111111;
				14'b01011100010111: oled_data = 16'b1111111111111111;
				14'b01011110010111: oled_data = 16'b1111111111111111;
				14'b01100000010111: oled_data = 16'b1111111111111111;
				14'b01100010010111: oled_data = 16'b1111111111111111;
				14'b01100100010111: oled_data = 16'b1111111111111111;
				14'b01100110010111: oled_data = 16'b1111111111111111;
				14'b01101000010111: oled_data = 16'b1111111111111111;
				14'b01101010010111: oled_data = 16'b1111111111111111;
				14'b01101100010111: oled_data = 16'b1111111111111111;
				14'b01101110010111: oled_data = 16'b1111111111111111;
				14'b01110000010111: oled_data = 16'b1111111111111111;
				14'b01110010010111: oled_data = 16'b1111111111111111;
				14'b01110100010111: oled_data = 16'b1111111111111111;
				14'b01110110010111: oled_data = 16'b1111111111111111;
				14'b01111000010111: oled_data = 16'b1111111111111111;
				14'b01111010010111: oled_data = 16'b1111111111111111;
				14'b01111100010111: oled_data = 16'b1111111111111111;
				14'b01111110010111: oled_data = 16'b1111111111111111;
				14'b10000000010111: oled_data = 16'b1111111111111111;
				14'b10000010010111: oled_data = 16'b1111111111111111;
				14'b10000100010111: oled_data = 16'b1111111111111111;
				14'b10000110010111: oled_data = 16'b1111111111111111;
				14'b10001000010111: oled_data = 16'b1111111111111111;
				14'b10001010010111: oled_data = 16'b1111111111111111;
				14'b10001100010111: oled_data = 16'b1111111111111111;
				14'b10001110010111: oled_data = 16'b1111111111111111;
				14'b10010000010111: oled_data = 16'b1111111111111111;
				14'b10010010010111: oled_data = 16'b1111111111111111;
				14'b10010100010111: oled_data = 16'b1111111111111111;
				14'b10010110010111: oled_data = 16'b1111111111111111;
				14'b10011000010111: oled_data = 16'b1111111111111111;
				14'b10011010010111: oled_data = 16'b1111111111111111;
				14'b10011100010111: oled_data = 16'b1111111111111111;
				14'b10011110010111: oled_data = 16'b1111111111111111;
				14'b10100000010111: oled_data = 16'b1111111111111111;
				14'b10100010010111: oled_data = 16'b1111111111111111;
				14'b10100100010111: oled_data = 16'b1111111111111111;
				14'b10100110010111: oled_data = 16'b1111111111111111;
				14'b10101000010111: oled_data = 16'b1111111111111111;
				14'b10101010010111: oled_data = 16'b1111111111111111;
				14'b10101100010111: oled_data = 16'b1111011111011110;
				14'b10101110010111: oled_data = 16'b1110011101111100;
				14'b10110000010111: oled_data = 16'b1100111100011001;
				14'b10110010010111: oled_data = 16'b1100111100011001;
				14'b10110100010111: oled_data = 16'b1101011100011001;
				14'b10110110010111: oled_data = 16'b1101011101011010;
				14'b10111000010111: oled_data = 16'b1101111101011011;
				14'b10111010010111: oled_data = 16'b1101111101011011;
				14'b10111100010111: oled_data = 16'b1101111101011011;
				14'b10111110010111: oled_data = 16'b1101111101011011;
				14'b00000000011000: oled_data = 16'b1111111111111111;
				14'b00000010011000: oled_data = 16'b1111111111111111;
				14'b00000100011000: oled_data = 16'b1111111111111111;
				14'b00000110011000: oled_data = 16'b1111111111111111;
				14'b00001000011000: oled_data = 16'b1111111111111111;
				14'b00001010011000: oled_data = 16'b1111111111111111;
				14'b00001100011000: oled_data = 16'b1111111111111111;
				14'b00001110011000: oled_data = 16'b1111111111111111;
				14'b00010000011000: oled_data = 16'b1111111111111111;
				14'b00010010011000: oled_data = 16'b1111111111111111;
				14'b00010100011000: oled_data = 16'b1111111111111111;
				14'b00010110011000: oled_data = 16'b1111111111111111;
				14'b00011000011000: oled_data = 16'b1111111111111111;
				14'b00011010011000: oled_data = 16'b1111111111111111;
				14'b00011100011000: oled_data = 16'b1111111111111111;
				14'b00011110011000: oled_data = 16'b1111111111111111;
				14'b00100000011000: oled_data = 16'b1111111111111111;
				14'b00100010011000: oled_data = 16'b1111111111111111;
				14'b00100100011000: oled_data = 16'b1111111111111111;
				14'b00100110011000: oled_data = 16'b1111111111111111;
				14'b00101000011000: oled_data = 16'b1111111111111111;
				14'b00101010011000: oled_data = 16'b1111111111111111;
				14'b00101100011000: oled_data = 16'b1111111111111111;
				14'b00101110011000: oled_data = 16'b1111111111111111;
				14'b00110000011000: oled_data = 16'b1111111111111111;
				14'b00110010011000: oled_data = 16'b1111111111111111;
				14'b00110100011000: oled_data = 16'b1111111111111111;
				14'b00110110011000: oled_data = 16'b1111111111111111;
				14'b00111000011000: oled_data = 16'b1111111111111111;
				14'b00111010011000: oled_data = 16'b1111111111111111;
				14'b00111100011000: oled_data = 16'b1111111111111111;
				14'b00111110011000: oled_data = 16'b1111111111111111;
				14'b01000000011000: oled_data = 16'b1111111111111111;
				14'b01000010011000: oled_data = 16'b1111111111111111;
				14'b01000100011000: oled_data = 16'b1111111111111111;
				14'b01000110011000: oled_data = 16'b1111111111111111;
				14'b01001000011000: oled_data = 16'b1111111111111111;
				14'b01001010011000: oled_data = 16'b1111111111111111;
				14'b01001100011000: oled_data = 16'b1111111111111111;
				14'b01001110011000: oled_data = 16'b1111111111111111;
				14'b01010000011000: oled_data = 16'b1111111111111111;
				14'b01010010011000: oled_data = 16'b1111111111111111;
				14'b01010100011000: oled_data = 16'b1111111111111111;
				14'b01010110011000: oled_data = 16'b1111111111111111;
				14'b01011000011000: oled_data = 16'b1111111111111111;
				14'b01011010011000: oled_data = 16'b1111111111111111;
				14'b01011100011000: oled_data = 16'b1111111111111111;
				14'b01011110011000: oled_data = 16'b1111111111111111;
				14'b01100000011000: oled_data = 16'b1111111111111111;
				14'b01100010011000: oled_data = 16'b1111111111111111;
				14'b01100100011000: oled_data = 16'b1111111111111111;
				14'b01100110011000: oled_data = 16'b1111111111111111;
				14'b01101000011000: oled_data = 16'b1111111111111111;
				14'b01101010011000: oled_data = 16'b1111111111111111;
				14'b01101100011000: oled_data = 16'b1111111111111111;
				14'b01101110011000: oled_data = 16'b1111111111111111;
				14'b01110000011000: oled_data = 16'b1111111111111111;
				14'b01110010011000: oled_data = 16'b1111111111111111;
				14'b01110100011000: oled_data = 16'b1111111111111111;
				14'b01110110011000: oled_data = 16'b1111111111111111;
				14'b01111000011000: oled_data = 16'b1111111111111111;
				14'b01111010011000: oled_data = 16'b1111111111111111;
				14'b01111100011000: oled_data = 16'b1111111111111111;
				14'b01111110011000: oled_data = 16'b1111111111111111;
				14'b10000000011000: oled_data = 16'b1111111111111111;
				14'b10000010011000: oled_data = 16'b1111111111111111;
				14'b10000100011000: oled_data = 16'b1111111111111111;
				14'b10000110011000: oled_data = 16'b1111111111111111;
				14'b10001000011000: oled_data = 16'b1111111111111111;
				14'b10001010011000: oled_data = 16'b1111111111111111;
				14'b10001100011000: oled_data = 16'b1111111111111111;
				14'b10001110011000: oled_data = 16'b1111111111111111;
				14'b10010000011000: oled_data = 16'b1111111111111111;
				14'b10010010011000: oled_data = 16'b1111111111111111;
				14'b10010100011000: oled_data = 16'b1111111111111111;
				14'b10010110011000: oled_data = 16'b1111111111111111;
				14'b10011000011000: oled_data = 16'b1111111111111111;
				14'b10011010011000: oled_data = 16'b1111111111111111;
				14'b10011100011000: oled_data = 16'b1111111111111111;
				14'b10011110011000: oled_data = 16'b1111111111111111;
				14'b10100000011000: oled_data = 16'b1111111111111111;
				14'b10100010011000: oled_data = 16'b1111111111111111;
				14'b10100100011000: oled_data = 16'b1111111111111111;
				14'b10100110011000: oled_data = 16'b1111111111111111;
				14'b10101000011000: oled_data = 16'b1111111111111111;
				14'b10101010011000: oled_data = 16'b1111111111111111;
				14'b10101100011000: oled_data = 16'b1111111111111111;
				14'b10101110011000: oled_data = 16'b1111011111011110;
				14'b10110000011000: oled_data = 16'b1110011110011100;
				14'b10110010011000: oled_data = 16'b1101011100111001;
				14'b10110100011000: oled_data = 16'b1100111100011000;
				14'b10110110011000: oled_data = 16'b1101011100011001;
				14'b10111000011000: oled_data = 16'b1101011100111010;
				14'b10111010011000: oled_data = 16'b1101111101011011;
				14'b10111100011000: oled_data = 16'b1101111101011011;
				14'b10111110011000: oled_data = 16'b1101111101011011;
				14'b00000000011001: oled_data = 16'b1111111111111111;
				14'b00000010011001: oled_data = 16'b1111111111111111;
				14'b00000100011001: oled_data = 16'b1111111111111111;
				14'b00000110011001: oled_data = 16'b1111111111111111;
				14'b00001000011001: oled_data = 16'b1111111111111111;
				14'b00001010011001: oled_data = 16'b1111111111111111;
				14'b00001100011001: oled_data = 16'b1111111111111111;
				14'b00001110011001: oled_data = 16'b1111111111111111;
				14'b00010000011001: oled_data = 16'b1111111111111111;
				14'b00010010011001: oled_data = 16'b1111111111111111;
				14'b00010100011001: oled_data = 16'b1111111111111111;
				14'b00010110011001: oled_data = 16'b1111111111111111;
				14'b00011000011001: oled_data = 16'b1111111111111111;
				14'b00011010011001: oled_data = 16'b1111111111111111;
				14'b00011100011001: oled_data = 16'b1111111111111111;
				14'b00011110011001: oled_data = 16'b1111111111111111;
				14'b00100000011001: oled_data = 16'b1111111111111111;
				14'b00100010011001: oled_data = 16'b1111111111111111;
				14'b00100100011001: oled_data = 16'b1111111111111111;
				14'b00100110011001: oled_data = 16'b1111111111111111;
				14'b00101000011001: oled_data = 16'b1111111111111111;
				14'b00101010011001: oled_data = 16'b1111111111111111;
				14'b00101100011001: oled_data = 16'b1111111111111111;
				14'b00101110011001: oled_data = 16'b1111111111111111;
				14'b00110000011001: oled_data = 16'b1111111111111111;
				14'b00110010011001: oled_data = 16'b1111111111111111;
				14'b00110100011001: oled_data = 16'b1111111111111111;
				14'b00110110011001: oled_data = 16'b1111111111111111;
				14'b00111000011001: oled_data = 16'b1111111111111111;
				14'b00111010011001: oled_data = 16'b1111111111111111;
				14'b00111100011001: oled_data = 16'b1111111111111111;
				14'b00111110011001: oled_data = 16'b1111111111111111;
				14'b01000000011001: oled_data = 16'b1111111111111111;
				14'b01000010011001: oled_data = 16'b1111111111111111;
				14'b01000100011001: oled_data = 16'b1111111111111111;
				14'b01000110011001: oled_data = 16'b1111111111111111;
				14'b01001000011001: oled_data = 16'b1111111111111111;
				14'b01001010011001: oled_data = 16'b1111111111111111;
				14'b01001100011001: oled_data = 16'b1111111111111111;
				14'b01001110011001: oled_data = 16'b1111111111111111;
				14'b01010000011001: oled_data = 16'b1111111111111111;
				14'b01010010011001: oled_data = 16'b1111111111111111;
				14'b01010100011001: oled_data = 16'b1111111111111111;
				14'b01010110011001: oled_data = 16'b1111111111111111;
				14'b01011000011001: oled_data = 16'b1111111111111111;
				14'b01011010011001: oled_data = 16'b1111111111111111;
				14'b01011100011001: oled_data = 16'b1111111111111111;
				14'b01011110011001: oled_data = 16'b1111111111111111;
				14'b01100000011001: oled_data = 16'b1111111111111111;
				14'b01100010011001: oled_data = 16'b1111111111111111;
				14'b01100100011001: oled_data = 16'b1111111111111111;
				14'b01100110011001: oled_data = 16'b1111111111111111;
				14'b01101000011001: oled_data = 16'b1111111111111111;
				14'b01101010011001: oled_data = 16'b1111111111111111;
				14'b01101100011001: oled_data = 16'b1111111111111111;
				14'b01101110011001: oled_data = 16'b1111111111111111;
				14'b01110000011001: oled_data = 16'b1111111111111111;
				14'b01110010011001: oled_data = 16'b1111111111111111;
				14'b01110100011001: oled_data = 16'b1111111111111111;
				14'b01110110011001: oled_data = 16'b1111111111111111;
				14'b01111000011001: oled_data = 16'b1111111111111111;
				14'b01111010011001: oled_data = 16'b1111111111111111;
				14'b01111100011001: oled_data = 16'b1111111111111111;
				14'b01111110011001: oled_data = 16'b1111111111111111;
				14'b10000000011001: oled_data = 16'b1111111111111111;
				14'b10000010011001: oled_data = 16'b1111111111111111;
				14'b10000100011001: oled_data = 16'b1111111111111111;
				14'b10000110011001: oled_data = 16'b1111111111111111;
				14'b10001000011001: oled_data = 16'b1111111111111111;
				14'b10001010011001: oled_data = 16'b1111111111111111;
				14'b10001100011001: oled_data = 16'b1111111111111111;
				14'b10001110011001: oled_data = 16'b1111111111111111;
				14'b10010000011001: oled_data = 16'b1111111111111111;
				14'b10010010011001: oled_data = 16'b1111111111111111;
				14'b10010100011001: oled_data = 16'b1111111111111111;
				14'b10010110011001: oled_data = 16'b1111111111111111;
				14'b10011000011001: oled_data = 16'b1111111111111111;
				14'b10011010011001: oled_data = 16'b1111111111111111;
				14'b10011100011001: oled_data = 16'b1111111111111111;
				14'b10011110011001: oled_data = 16'b1111111111111111;
				14'b10100000011001: oled_data = 16'b1111111111111111;
				14'b10100010011001: oled_data = 16'b1111111111111111;
				14'b10100100011001: oled_data = 16'b1111111111111111;
				14'b10100110011001: oled_data = 16'b1111111111111111;
				14'b10101000011001: oled_data = 16'b1111111111111111;
				14'b10101010011001: oled_data = 16'b1111111111111111;
				14'b10101100011001: oled_data = 16'b1111111111111111;
				14'b10101110011001: oled_data = 16'b1111111111111111;
				14'b10110000011001: oled_data = 16'b1111111111111111;
				14'b10110010011001: oled_data = 16'b1110111110111101;
				14'b10110100011001: oled_data = 16'b1101011100111010;
				14'b10110110011001: oled_data = 16'b1100111100011000;
				14'b10111000011001: oled_data = 16'b1101011100011001;
				14'b10111010011001: oled_data = 16'b1101011100111001;
				14'b10111100011001: oled_data = 16'b1101111101011010;
				14'b10111110011001: oled_data = 16'b1101111101011011;
				14'b00000000011010: oled_data = 16'b1111111111111111;
				14'b00000010011010: oled_data = 16'b1111111111111111;
				14'b00000100011010: oled_data = 16'b1111111111111111;
				14'b00000110011010: oled_data = 16'b1111111111111111;
				14'b00001000011010: oled_data = 16'b1111111111111111;
				14'b00001010011010: oled_data = 16'b1111111111111111;
				14'b00001100011010: oled_data = 16'b1111111111111111;
				14'b00001110011010: oled_data = 16'b1111111111111111;
				14'b00010000011010: oled_data = 16'b1111111111111111;
				14'b00010010011010: oled_data = 16'b1111111111111111;
				14'b00010100011010: oled_data = 16'b1111111111111111;
				14'b00010110011010: oled_data = 16'b1111111111111111;
				14'b00011000011010: oled_data = 16'b1111111111111111;
				14'b00011010011010: oled_data = 16'b1111111111111111;
				14'b00011100011010: oled_data = 16'b1111111111111111;
				14'b00011110011010: oled_data = 16'b1111111111111111;
				14'b00100000011010: oled_data = 16'b1111111111111111;
				14'b00100010011010: oled_data = 16'b1111111111111111;
				14'b00100100011010: oled_data = 16'b1111111111111111;
				14'b00100110011010: oled_data = 16'b1111111111111111;
				14'b00101000011010: oled_data = 16'b1111111111111111;
				14'b00101010011010: oled_data = 16'b1111111111111111;
				14'b00101100011010: oled_data = 16'b1111111111111111;
				14'b00101110011010: oled_data = 16'b1111111111111111;
				14'b00110000011010: oled_data = 16'b1111111111111111;
				14'b00110010011010: oled_data = 16'b1111111111111111;
				14'b00110100011010: oled_data = 16'b1111111111111111;
				14'b00110110011010: oled_data = 16'b1111111111111111;
				14'b00111000011010: oled_data = 16'b1111111111111111;
				14'b00111010011010: oled_data = 16'b1111111111111111;
				14'b00111100011010: oled_data = 16'b1111111111111111;
				14'b00111110011010: oled_data = 16'b1111111111111111;
				14'b01000000011010: oled_data = 16'b1111111111111111;
				14'b01000010011010: oled_data = 16'b1111111111111111;
				14'b01000100011010: oled_data = 16'b1111111111111111;
				14'b01000110011010: oled_data = 16'b1111111111111111;
				14'b01001000011010: oled_data = 16'b1111111111111111;
				14'b01001010011010: oled_data = 16'b1111111111111111;
				14'b01001100011010: oled_data = 16'b1111111111111111;
				14'b01001110011010: oled_data = 16'b1111111111111111;
				14'b01010000011010: oled_data = 16'b1111111111111111;
				14'b01010010011010: oled_data = 16'b1111111111111111;
				14'b01010100011010: oled_data = 16'b1111111111111111;
				14'b01010110011010: oled_data = 16'b1111111111111111;
				14'b01011000011010: oled_data = 16'b1111111111111111;
				14'b01011010011010: oled_data = 16'b1111111111111111;
				14'b01011100011010: oled_data = 16'b1111111111111111;
				14'b01011110011010: oled_data = 16'b1111111111111111;
				14'b01100000011010: oled_data = 16'b1111111111111111;
				14'b01100010011010: oled_data = 16'b1111111111111111;
				14'b01100100011010: oled_data = 16'b1111111111111111;
				14'b01100110011010: oled_data = 16'b1111111111111111;
				14'b01101000011010: oled_data = 16'b1111111111111111;
				14'b01101010011010: oled_data = 16'b1111111111111111;
				14'b01101100011010: oled_data = 16'b1111111111111111;
				14'b01101110011010: oled_data = 16'b1111111111111111;
				14'b01110000011010: oled_data = 16'b1111111111111111;
				14'b01110010011010: oled_data = 16'b1111111111111111;
				14'b01110100011010: oled_data = 16'b1111111111111111;
				14'b01110110011010: oled_data = 16'b1111111111111111;
				14'b01111000011010: oled_data = 16'b1111111111111111;
				14'b01111010011010: oled_data = 16'b1111111111111111;
				14'b01111100011010: oled_data = 16'b1111111111111111;
				14'b01111110011010: oled_data = 16'b1111111111111111;
				14'b10000000011010: oled_data = 16'b1111111111111111;
				14'b10000010011010: oled_data = 16'b1111111111111111;
				14'b10000100011010: oled_data = 16'b1111111111111111;
				14'b10000110011010: oled_data = 16'b1111111111111111;
				14'b10001000011010: oled_data = 16'b1111111111111111;
				14'b10001010011010: oled_data = 16'b1111111111111111;
				14'b10001100011010: oled_data = 16'b1111111111111111;
				14'b10001110011010: oled_data = 16'b1111111111111111;
				14'b10010000011010: oled_data = 16'b1111111111111111;
				14'b10010010011010: oled_data = 16'b1111111111111111;
				14'b10010100011010: oled_data = 16'b1111111111111111;
				14'b10010110011010: oled_data = 16'b1111111111111111;
				14'b10011000011010: oled_data = 16'b1111111111111111;
				14'b10011010011010: oled_data = 16'b1111111111111111;
				14'b10011100011010: oled_data = 16'b1111111111111111;
				14'b10011110011010: oled_data = 16'b1111111111111111;
				14'b10100000011010: oled_data = 16'b1111111111111111;
				14'b10100010011010: oled_data = 16'b1111111111111111;
				14'b10100100011010: oled_data = 16'b1111111111111111;
				14'b10100110011010: oled_data = 16'b1111111111111111;
				14'b10101000011010: oled_data = 16'b1111111111111111;
				14'b10101010011010: oled_data = 16'b1111111111111111;
				14'b10101100011010: oled_data = 16'b1111111111111111;
				14'b10101110011010: oled_data = 16'b1111111111111111;
				14'b10110000011010: oled_data = 16'b1111111111111111;
				14'b10110010011010: oled_data = 16'b1111111111111111;
				14'b10110100011010: oled_data = 16'b1111011111011110;
				14'b10110110011010: oled_data = 16'b1110011101111011;
				14'b10111000011010: oled_data = 16'b1101011100011001;
				14'b10111010011010: oled_data = 16'b1100111100011000;
				14'b10111100011010: oled_data = 16'b1101011100111001;
				14'b10111110011010: oled_data = 16'b1101011100111001;
				14'b00000000011011: oled_data = 16'b1111111111111111;
				14'b00000010011011: oled_data = 16'b1111111111111111;
				14'b00000100011011: oled_data = 16'b1111111111111111;
				14'b00000110011011: oled_data = 16'b1111111111111111;
				14'b00001000011011: oled_data = 16'b1111111111111111;
				14'b00001010011011: oled_data = 16'b1111111111111111;
				14'b00001100011011: oled_data = 16'b1111111111111111;
				14'b00001110011011: oled_data = 16'b1111111111111111;
				14'b00010000011011: oled_data = 16'b1111111111111111;
				14'b00010010011011: oled_data = 16'b1111111111111111;
				14'b00010100011011: oled_data = 16'b1111111111111111;
				14'b00010110011011: oled_data = 16'b1111111111111111;
				14'b00011000011011: oled_data = 16'b1111111111111111;
				14'b00011010011011: oled_data = 16'b1111111111111111;
				14'b00011100011011: oled_data = 16'b1111111111111111;
				14'b00011110011011: oled_data = 16'b1111111111111111;
				14'b00100000011011: oled_data = 16'b1111111111111111;
				14'b00100010011011: oled_data = 16'b1111111111111111;
				14'b00100100011011: oled_data = 16'b1111111111111111;
				14'b00100110011011: oled_data = 16'b1111111111111111;
				14'b00101000011011: oled_data = 16'b1111111111111111;
				14'b00101010011011: oled_data = 16'b1111111111111111;
				14'b00101100011011: oled_data = 16'b1111111111111111;
				14'b00101110011011: oled_data = 16'b1111111111111111;
				14'b00110000011011: oled_data = 16'b1111111111111111;
				14'b00110010011011: oled_data = 16'b1111111111111111;
				14'b00110100011011: oled_data = 16'b1111111111111111;
				14'b00110110011011: oled_data = 16'b1111111111111111;
				14'b00111000011011: oled_data = 16'b1111111111111111;
				14'b00111010011011: oled_data = 16'b1111111111111111;
				14'b00111100011011: oled_data = 16'b1111111111111111;
				14'b00111110011011: oled_data = 16'b1111111111111111;
				14'b01000000011011: oled_data = 16'b1111111111111111;
				14'b01000010011011: oled_data = 16'b1111111111111111;
				14'b01000100011011: oled_data = 16'b1111111111111111;
				14'b01000110011011: oled_data = 16'b1111111111111111;
				14'b01001000011011: oled_data = 16'b1111111111111111;
				14'b01001010011011: oled_data = 16'b1111111111111111;
				14'b01001100011011: oled_data = 16'b1111111111111111;
				14'b01001110011011: oled_data = 16'b1111111111111111;
				14'b01010000011011: oled_data = 16'b1111111111111111;
				14'b01010010011011: oled_data = 16'b1111111111111111;
				14'b01010100011011: oled_data = 16'b1111111111111111;
				14'b01010110011011: oled_data = 16'b1111111111111111;
				14'b01011000011011: oled_data = 16'b1111111111111111;
				14'b01011010011011: oled_data = 16'b1111111111111111;
				14'b01011100011011: oled_data = 16'b1111111111111111;
				14'b01011110011011: oled_data = 16'b1111111111111111;
				14'b01100000011011: oled_data = 16'b1111111111111111;
				14'b01100010011011: oled_data = 16'b1111111111111111;
				14'b01100100011011: oled_data = 16'b1111111111111111;
				14'b01100110011011: oled_data = 16'b1111111111111111;
				14'b01101000011011: oled_data = 16'b1111111111111111;
				14'b01101010011011: oled_data = 16'b1111111111111111;
				14'b01101100011011: oled_data = 16'b1111111111111111;
				14'b01101110011011: oled_data = 16'b1111111111111111;
				14'b01110000011011: oled_data = 16'b1111111111111111;
				14'b01110010011011: oled_data = 16'b1111111111111111;
				14'b01110100011011: oled_data = 16'b1111111111111111;
				14'b01110110011011: oled_data = 16'b1111111111111111;
				14'b01111000011011: oled_data = 16'b1111111111111111;
				14'b01111010011011: oled_data = 16'b1111111111111111;
				14'b01111100011011: oled_data = 16'b1111111111111111;
				14'b01111110011011: oled_data = 16'b1111111111111111;
				14'b10000000011011: oled_data = 16'b1111111111111111;
				14'b10000010011011: oled_data = 16'b1111111111111111;
				14'b10000100011011: oled_data = 16'b1111111111111111;
				14'b10000110011011: oled_data = 16'b1111111111111111;
				14'b10001000011011: oled_data = 16'b1111111111111111;
				14'b10001010011011: oled_data = 16'b1111111111111111;
				14'b10001100011011: oled_data = 16'b1111111111111111;
				14'b10001110011011: oled_data = 16'b1111111111111111;
				14'b10010000011011: oled_data = 16'b1111111111111111;
				14'b10010010011011: oled_data = 16'b1111111111111111;
				14'b10010100011011: oled_data = 16'b1111111111111111;
				14'b10010110011011: oled_data = 16'b1111111111111111;
				14'b10011000011011: oled_data = 16'b1111111111111111;
				14'b10011010011011: oled_data = 16'b1111111111111111;
				14'b10011100011011: oled_data = 16'b1111111111111111;
				14'b10011110011011: oled_data = 16'b1111111111111111;
				14'b10100000011011: oled_data = 16'b1111111111111111;
				14'b10100010011011: oled_data = 16'b1111111111111111;
				14'b10100100011011: oled_data = 16'b1111111111111111;
				14'b10100110011011: oled_data = 16'b1111111111111111;
				14'b10101000011011: oled_data = 16'b1111111111111111;
				14'b10101010011011: oled_data = 16'b1111111111111111;
				14'b10101100011011: oled_data = 16'b1111111111111111;
				14'b10101110011011: oled_data = 16'b1111111111111111;
				14'b10110000011011: oled_data = 16'b1111111111111111;
				14'b10110010011011: oled_data = 16'b1111111111111111;
				14'b10110100011011: oled_data = 16'b1111111111111111;
				14'b10110110011011: oled_data = 16'b1111111111111111;
				14'b10111000011011: oled_data = 16'b1111011111011110;
				14'b10111010011011: oled_data = 16'b1101111101111011;
				14'b10111100011011: oled_data = 16'b1101011100111001;
				14'b10111110011011: oled_data = 16'b1100111100011000;
				14'b00000000011100: oled_data = 16'b1111111111111111;
				14'b00000010011100: oled_data = 16'b1111111111111111;
				14'b00000100011100: oled_data = 16'b1111111111111111;
				14'b00000110011100: oled_data = 16'b1111111111111111;
				14'b00001000011100: oled_data = 16'b1111111111111111;
				14'b00001010011100: oled_data = 16'b1111111111111111;
				14'b00001100011100: oled_data = 16'b1111111111111111;
				14'b00001110011100: oled_data = 16'b1111111111111111;
				14'b00010000011100: oled_data = 16'b1111111111111111;
				14'b00010010011100: oled_data = 16'b1111111111111111;
				14'b00010100011100: oled_data = 16'b1111111111111111;
				14'b00010110011100: oled_data = 16'b1111111111111111;
				14'b00011000011100: oled_data = 16'b1111111111111111;
				14'b00011010011100: oled_data = 16'b1111111111111111;
				14'b00011100011100: oled_data = 16'b1111111111111111;
				14'b00011110011100: oled_data = 16'b1111111111111111;
				14'b00100000011100: oled_data = 16'b1111111111111111;
				14'b00100010011100: oled_data = 16'b1111111111111111;
				14'b00100100011100: oled_data = 16'b1111111111111111;
				14'b00100110011100: oled_data = 16'b1111111111111111;
				14'b00101000011100: oled_data = 16'b1111111111111111;
				14'b00101010011100: oled_data = 16'b1111111111111111;
				14'b00101100011100: oled_data = 16'b1111111111111111;
				14'b00101110011100: oled_data = 16'b1111111111111111;
				14'b00110000011100: oled_data = 16'b1111111111111111;
				14'b00110010011100: oled_data = 16'b1111111111111111;
				14'b00110100011100: oled_data = 16'b1111111111111111;
				14'b00110110011100: oled_data = 16'b1111111111111111;
				14'b00111000011100: oled_data = 16'b1111111111111111;
				14'b00111010011100: oled_data = 16'b1111111111111111;
				14'b00111100011100: oled_data = 16'b1111111111111111;
				14'b00111110011100: oled_data = 16'b1111111111111111;
				14'b01000000011100: oled_data = 16'b1111111111111111;
				14'b01000010011100: oled_data = 16'b1111111111111111;
				14'b01000100011100: oled_data = 16'b1111111111111111;
				14'b01000110011100: oled_data = 16'b1111111111111111;
				14'b01001000011100: oled_data = 16'b1111111111111111;
				14'b01001010011100: oled_data = 16'b1111111111111111;
				14'b01001100011100: oled_data = 16'b1111111111111111;
				14'b01001110011100: oled_data = 16'b1111111111111111;
				14'b01010000011100: oled_data = 16'b1111111111111111;
				14'b01010010011100: oled_data = 16'b1111111111111111;
				14'b01010100011100: oled_data = 16'b1111111111111111;
				14'b01010110011100: oled_data = 16'b1111111111111111;
				14'b01011000011100: oled_data = 16'b1111111111111111;
				14'b01011010011100: oled_data = 16'b1111111111111111;
				14'b01011100011100: oled_data = 16'b1111111111111111;
				14'b01011110011100: oled_data = 16'b1111111111111111;
				14'b01100000011100: oled_data = 16'b1111111111111111;
				14'b01100010011100: oled_data = 16'b1111111111111111;
				14'b01100100011100: oled_data = 16'b1111111111111111;
				14'b01100110011100: oled_data = 16'b1111111111111111;
				14'b01101000011100: oled_data = 16'b1111111111111111;
				14'b01101010011100: oled_data = 16'b1111111111111111;
				14'b01101100011100: oled_data = 16'b1111111111111111;
				14'b01101110011100: oled_data = 16'b1111111111111111;
				14'b01110000011100: oled_data = 16'b1111111111111111;
				14'b01110010011100: oled_data = 16'b1111111111111111;
				14'b01110100011100: oled_data = 16'b1111111111111111;
				14'b01110110011100: oled_data = 16'b1111111111111111;
				14'b01111000011100: oled_data = 16'b1111111111111111;
				14'b01111010011100: oled_data = 16'b1111111111111111;
				14'b01111100011100: oled_data = 16'b1111111111111111;
				14'b01111110011100: oled_data = 16'b1111111111111111;
				14'b10000000011100: oled_data = 16'b1111111111111111;
				14'b10000010011100: oled_data = 16'b1111111111111111;
				14'b10000100011100: oled_data = 16'b1111111111111111;
				14'b10000110011100: oled_data = 16'b1111111111111111;
				14'b10001000011100: oled_data = 16'b1111111111111111;
				14'b10001010011100: oled_data = 16'b1111111111111111;
				14'b10001100011100: oled_data = 16'b1111111111111111;
				14'b10001110011100: oled_data = 16'b1111111111111111;
				14'b10010000011100: oled_data = 16'b1111111111111111;
				14'b10010010011100: oled_data = 16'b1111111111111111;
				14'b10010100011100: oled_data = 16'b1111111111111111;
				14'b10010110011100: oled_data = 16'b1111111111111111;
				14'b10011000011100: oled_data = 16'b1111111111111111;
				14'b10011010011100: oled_data = 16'b1111111111111111;
				14'b10011100011100: oled_data = 16'b1111111111111111;
				14'b10011110011100: oled_data = 16'b1111111111111111;
				14'b10100000011100: oled_data = 16'b1111111111111111;
				14'b10100010011100: oled_data = 16'b1111111111111111;
				14'b10100100011100: oled_data = 16'b1111111111111111;
				14'b10100110011100: oled_data = 16'b1111111111111111;
				14'b10101000011100: oled_data = 16'b1111111111111111;
				14'b10101010011100: oled_data = 16'b1111111111111111;
				14'b10101100011100: oled_data = 16'b1111111111111111;
				14'b10101110011100: oled_data = 16'b1111111111111111;
				14'b10110000011100: oled_data = 16'b1111111111111111;
				14'b10110010011100: oled_data = 16'b1111111111111111;
				14'b10110100011100: oled_data = 16'b1111111111111111;
				14'b10110110011100: oled_data = 16'b1111111111111111;
				14'b10111000011100: oled_data = 16'b1111111111111111;
				14'b10111010011100: oled_data = 16'b1111111111111111;
				14'b10111100011100: oled_data = 16'b1111011111011110;
				14'b10111110011100: oled_data = 16'b1110111110011100;
				14'b00000000011101: oled_data = 16'b1111111111111111;
				14'b00000010011101: oled_data = 16'b1111111111111111;
				14'b00000100011101: oled_data = 16'b1111111111111111;
				14'b00000110011101: oled_data = 16'b1111111111111111;
				14'b00001000011101: oled_data = 16'b1111111111111111;
				14'b00001010011101: oled_data = 16'b1111111111111111;
				14'b00001100011101: oled_data = 16'b1111111111111111;
				14'b00001110011101: oled_data = 16'b1111111111111111;
				14'b00010000011101: oled_data = 16'b1111111111111111;
				14'b00010010011101: oled_data = 16'b1111111111111111;
				14'b00010100011101: oled_data = 16'b1111111111111111;
				14'b00010110011101: oled_data = 16'b1111111111111111;
				14'b00011000011101: oled_data = 16'b1111111111111111;
				14'b00011010011101: oled_data = 16'b1111111111111111;
				14'b00011100011101: oled_data = 16'b1111111111111111;
				14'b00011110011101: oled_data = 16'b1111111111111111;
				14'b00100000011101: oled_data = 16'b1111111111111111;
				14'b00100010011101: oled_data = 16'b1111111111111111;
				14'b00100100011101: oled_data = 16'b1111111111111111;
				14'b00100110011101: oled_data = 16'b1111111111111111;
				14'b00101000011101: oled_data = 16'b1111111111111111;
				14'b00101010011101: oled_data = 16'b1111111111111111;
				14'b00101100011101: oled_data = 16'b1111111111111111;
				14'b00101110011101: oled_data = 16'b1111111111111111;
				14'b00110000011101: oled_data = 16'b1111111111111111;
				14'b00110010011101: oled_data = 16'b1111111111111111;
				14'b00110100011101: oled_data = 16'b1111111111111111;
				14'b00110110011101: oled_data = 16'b1111111111111111;
				14'b00111000011101: oled_data = 16'b1111111111111111;
				14'b00111010011101: oled_data = 16'b1111111111111111;
				14'b00111100011101: oled_data = 16'b1111111111111111;
				14'b00111110011101: oled_data = 16'b1111111111111111;
				14'b01000000011101: oled_data = 16'b1111111111111111;
				14'b01000010011101: oled_data = 16'b1111111111111111;
				14'b01000100011101: oled_data = 16'b1111111111111111;
				14'b01000110011101: oled_data = 16'b1111111111111111;
				14'b01001000011101: oled_data = 16'b1111111111111111;
				14'b01001010011101: oled_data = 16'b1111111111111111;
				14'b01001100011101: oled_data = 16'b1111111111111111;
				14'b01001110011101: oled_data = 16'b1111111111111111;
				14'b01010000011101: oled_data = 16'b1111111111111111;
				14'b01010010011101: oled_data = 16'b1111111111111111;
				14'b01010100011101: oled_data = 16'b1111111111111111;
				14'b01010110011101: oled_data = 16'b1111111111111111;
				14'b01011000011101: oled_data = 16'b1111111111111111;
				14'b01011010011101: oled_data = 16'b1111111111111111;
				14'b01011100011101: oled_data = 16'b1111111111111111;
				14'b01011110011101: oled_data = 16'b1111111111111111;
				14'b01100000011101: oled_data = 16'b1111111111111111;
				14'b01100010011101: oled_data = 16'b1111111111111111;
				14'b01100100011101: oled_data = 16'b1111111111111111;
				14'b01100110011101: oled_data = 16'b1111111111111111;
				14'b01101000011101: oled_data = 16'b1111111111111111;
				14'b01101010011101: oled_data = 16'b1111111111111111;
				14'b01101100011101: oled_data = 16'b1111111111111111;
				14'b01101110011101: oled_data = 16'b1111111111111111;
				14'b01110000011101: oled_data = 16'b1111111111111111;
				14'b01110010011101: oled_data = 16'b1111111111111111;
				14'b01110100011101: oled_data = 16'b1111111111111111;
				14'b01110110011101: oled_data = 16'b1111111111111111;
				14'b01111000011101: oled_data = 16'b1111111111111111;
				14'b01111010011101: oled_data = 16'b1111111111111111;
				14'b01111100011101: oled_data = 16'b1111111111111111;
				14'b01111110011101: oled_data = 16'b1111111111111111;
				14'b10000000011101: oled_data = 16'b1111111111111111;
				14'b10000010011101: oled_data = 16'b1111111111111111;
				14'b10000100011101: oled_data = 16'b1111111111111111;
				14'b10000110011101: oled_data = 16'b1111111111111111;
				14'b10001000011101: oled_data = 16'b1111111111111111;
				14'b10001010011101: oled_data = 16'b1111111111111111;
				14'b10001100011101: oled_data = 16'b1111111111111111;
				14'b10001110011101: oled_data = 16'b1111111111111111;
				14'b10010000011101: oled_data = 16'b1111111111111111;
				14'b10010010011101: oled_data = 16'b1111111111111111;
				14'b10010100011101: oled_data = 16'b1111111111111111;
				14'b10010110011101: oled_data = 16'b1111111111111111;
				14'b10011000011101: oled_data = 16'b1111111111111111;
				14'b10011010011101: oled_data = 16'b1111111111111111;
				14'b10011100011101: oled_data = 16'b1111111111111111;
				14'b10011110011101: oled_data = 16'b1111111111111111;
				14'b10100000011101: oled_data = 16'b1111111111111111;
				14'b10100010011101: oled_data = 16'b1111111111111111;
				14'b10100100011101: oled_data = 16'b1111111111111111;
				14'b10100110011101: oled_data = 16'b1111111111111111;
				14'b10101000011101: oled_data = 16'b1111111111111111;
				14'b10101010011101: oled_data = 16'b1111111111111111;
				14'b10101100011101: oled_data = 16'b1111111111111111;
				14'b10101110011101: oled_data = 16'b1111111111111111;
				14'b10110000011101: oled_data = 16'b1111111111111111;
				14'b10110010011101: oled_data = 16'b1111111111111111;
				14'b10110100011101: oled_data = 16'b1111111111111111;
				14'b10110110011101: oled_data = 16'b1111111111111111;
				14'b10111000011101: oled_data = 16'b1111111111111111;
				14'b10111010011101: oled_data = 16'b1111111111111111;
				14'b10111100011101: oled_data = 16'b1111111111111111;
				14'b10111110011101: oled_data = 16'b1111111111111111;
				14'b00000000011110: oled_data = 16'b1111111111111111;
				14'b00000010011110: oled_data = 16'b1111111111111111;
				14'b00000100011110: oled_data = 16'b1111111111111111;
				14'b00000110011110: oled_data = 16'b1111111111111111;
				14'b00001000011110: oled_data = 16'b1111111111111111;
				14'b00001010011110: oled_data = 16'b1111111111111111;
				14'b00001100011110: oled_data = 16'b1111111111111111;
				14'b00001110011110: oled_data = 16'b1111111111111111;
				14'b00010000011110: oled_data = 16'b1111111111111111;
				14'b00010010011110: oled_data = 16'b1111111111111111;
				14'b00010100011110: oled_data = 16'b1111111111111111;
				14'b00010110011110: oled_data = 16'b1111111111111111;
				14'b00011000011110: oled_data = 16'b1111111111111111;
				14'b00011010011110: oled_data = 16'b1111111111111111;
				14'b00011100011110: oled_data = 16'b1111111111111111;
				14'b00011110011110: oled_data = 16'b1111111111111111;
				14'b00100000011110: oled_data = 16'b1111111111111111;
				14'b00100010011110: oled_data = 16'b1111111111111111;
				14'b00100100011110: oled_data = 16'b1111111111111111;
				14'b00100110011110: oled_data = 16'b1111111111111111;
				14'b00101000011110: oled_data = 16'b1111111111111111;
				14'b00101010011110: oled_data = 16'b1111111111111111;
				14'b00101100011110: oled_data = 16'b1111111111111111;
				14'b00101110011110: oled_data = 16'b1111111111111111;
				14'b00110000011110: oled_data = 16'b1111111111111111;
				14'b00110010011110: oled_data = 16'b1111111111111111;
				14'b00110100011110: oled_data = 16'b1111111111111111;
				14'b00110110011110: oled_data = 16'b1111111111111111;
				14'b00111000011110: oled_data = 16'b1111111111111111;
				14'b00111010011110: oled_data = 16'b1111111111111111;
				14'b00111100011110: oled_data = 16'b1111111111111111;
				14'b00111110011110: oled_data = 16'b1111111111111111;
				14'b01000000011110: oled_data = 16'b1111111111111111;
				14'b01000010011110: oled_data = 16'b1111111111111111;
				14'b01000100011110: oled_data = 16'b1111111111111111;
				14'b01000110011110: oled_data = 16'b1111111111111111;
				14'b01001000011110: oled_data = 16'b1111111111111111;
				14'b01001010011110: oled_data = 16'b1111111111111111;
				14'b01001100011110: oled_data = 16'b1111111111111111;
				14'b01001110011110: oled_data = 16'b1111111111111111;
				14'b01010000011110: oled_data = 16'b1111111111111111;
				14'b01010010011110: oled_data = 16'b1111111111111111;
				14'b01010100011110: oled_data = 16'b1111111111111111;
				14'b01010110011110: oled_data = 16'b1111111111111111;
				14'b01011000011110: oled_data = 16'b1111111111111111;
				14'b01011010011110: oled_data = 16'b1111111111111111;
				14'b01011100011110: oled_data = 16'b1111111111111111;
				14'b01011110011110: oled_data = 16'b1111111111111111;
				14'b01100000011110: oled_data = 16'b1111111111111111;
				14'b01100010011110: oled_data = 16'b1111111111111111;
				14'b01100100011110: oled_data = 16'b1111111111111111;
				14'b01100110011110: oled_data = 16'b1111111111111111;
				14'b01101000011110: oled_data = 16'b1111111111111111;
				14'b01101010011110: oled_data = 16'b1111111111111111;
				14'b01101100011110: oled_data = 16'b1111111111111111;
				14'b01101110011110: oled_data = 16'b1111111111111111;
				14'b01110000011110: oled_data = 16'b1111111111111111;
				14'b01110010011110: oled_data = 16'b1111111111111111;
				14'b01110100011110: oled_data = 16'b1111111111111111;
				14'b01110110011110: oled_data = 16'b1111111111111111;
				14'b01111000011110: oled_data = 16'b1111111111111111;
				14'b01111010011110: oled_data = 16'b1111111111111111;
				14'b01111100011110: oled_data = 16'b1111111111111111;
				14'b01111110011110: oled_data = 16'b1111111111111111;
				14'b10000000011110: oled_data = 16'b1111111111111111;
				14'b10000010011110: oled_data = 16'b1111111111111111;
				14'b10000100011110: oled_data = 16'b1111111111111111;
				14'b10000110011110: oled_data = 16'b1111111111111111;
				14'b10001000011110: oled_data = 16'b1111111111111111;
				14'b10001010011110: oled_data = 16'b1111111111111111;
				14'b10001100011110: oled_data = 16'b1111111111111111;
				14'b10001110011110: oled_data = 16'b1111111111111111;
				14'b10010000011110: oled_data = 16'b1111111111111111;
				14'b10010010011110: oled_data = 16'b1111111111111111;
				14'b10010100011110: oled_data = 16'b1111111111111111;
				14'b10010110011110: oled_data = 16'b1111111111111111;
				14'b10011000011110: oled_data = 16'b1111111111111111;
				14'b10011010011110: oled_data = 16'b1111111111111111;
				14'b10011100011110: oled_data = 16'b1111111111111111;
				14'b10011110011110: oled_data = 16'b1111111111111111;
				14'b10100000011110: oled_data = 16'b1111111111111111;
				14'b10100010011110: oled_data = 16'b1111111111111111;
				14'b10100100011110: oled_data = 16'b1111111111111111;
				14'b10100110011110: oled_data = 16'b1111111111111111;
				14'b10101000011110: oled_data = 16'b1111111111111111;
				14'b10101010011110: oled_data = 16'b1111111111111111;
				14'b10101100011110: oled_data = 16'b1111111111111111;
				14'b10101110011110: oled_data = 16'b1111111111111111;
				14'b10110000011110: oled_data = 16'b1111111111111111;
				14'b10110010011110: oled_data = 16'b1111111111111111;
				14'b10110100011110: oled_data = 16'b1111111111111111;
				14'b10110110011110: oled_data = 16'b1111111111111111;
				14'b10111000011110: oled_data = 16'b1111111111111111;
				14'b10111010011110: oled_data = 16'b1111111111111111;
				14'b10111100011110: oled_data = 16'b1111111111111111;
				14'b10111110011110: oled_data = 16'b1111111111111111;
				14'b00000000011111: oled_data = 16'b1111111111111111;
				14'b00000010011111: oled_data = 16'b1111111111111111;
				14'b00000100011111: oled_data = 16'b1111111111111111;
				14'b00000110011111: oled_data = 16'b1111111111111111;
				14'b00001000011111: oled_data = 16'b1111111111111111;
				14'b00001010011111: oled_data = 16'b1111111111111111;
				14'b00001100011111: oled_data = 16'b1111111111111111;
				14'b00001110011111: oled_data = 16'b1111111111111111;
				14'b00010000011111: oled_data = 16'b1111111111111111;
				14'b00010010011111: oled_data = 16'b1111111111111111;
				14'b00010100011111: oled_data = 16'b1111111111111111;
				14'b00010110011111: oled_data = 16'b1111111111111111;
				14'b00011000011111: oled_data = 16'b1111111111111111;
				14'b00011010011111: oled_data = 16'b1111111111111111;
				14'b00011100011111: oled_data = 16'b1111111111111111;
				14'b00011110011111: oled_data = 16'b1111111111111111;
				14'b00100000011111: oled_data = 16'b1111111111111111;
				14'b00100010011111: oled_data = 16'b1111111111111111;
				14'b00100100011111: oled_data = 16'b1111111111111111;
				14'b00100110011111: oled_data = 16'b1111111111111111;
				14'b00101000011111: oled_data = 16'b1111111111111111;
				14'b00101010011111: oled_data = 16'b1111111111111111;
				14'b00101100011111: oled_data = 16'b1111111111111111;
				14'b00101110011111: oled_data = 16'b1111111111111111;
				14'b00110000011111: oled_data = 16'b1111111111111111;
				14'b00110010011111: oled_data = 16'b1111111111111111;
				14'b00110100011111: oled_data = 16'b1111111111111111;
				14'b00110110011111: oled_data = 16'b1111111111111111;
				14'b00111000011111: oled_data = 16'b1111111111111111;
				14'b00111010011111: oled_data = 16'b1111111111111111;
				14'b00111100011111: oled_data = 16'b1111111111111111;
				14'b00111110011111: oled_data = 16'b1111111111111111;
				14'b01000000011111: oled_data = 16'b1111111111111111;
				14'b01000010011111: oled_data = 16'b1111111111111111;
				14'b01000100011111: oled_data = 16'b1111111111111111;
				14'b01000110011111: oled_data = 16'b1111111111111111;
				14'b01001000011111: oled_data = 16'b1111111111111111;
				14'b01001010011111: oled_data = 16'b1111111111111111;
				14'b01001100011111: oled_data = 16'b1111111111111111;
				14'b01001110011111: oled_data = 16'b1111111111111111;
				14'b01010000011111: oled_data = 16'b1111111111111111;
				14'b01010010011111: oled_data = 16'b1111111111111111;
				14'b01010100011111: oled_data = 16'b1111111111111111;
				14'b01010110011111: oled_data = 16'b1111111111111111;
				14'b01011000011111: oled_data = 16'b1111111111111111;
				14'b01011010011111: oled_data = 16'b1111111111111111;
				14'b01011100011111: oled_data = 16'b1111111111111111;
				14'b01011110011111: oled_data = 16'b1111111111111111;
				14'b01100000011111: oled_data = 16'b1111111111111111;
				14'b01100010011111: oled_data = 16'b1111111111111111;
				14'b01100100011111: oled_data = 16'b1111111111111111;
				14'b01100110011111: oled_data = 16'b1111111111111111;
				14'b01101000011111: oled_data = 16'b1111111111111111;
				14'b01101010011111: oled_data = 16'b1111111111111111;
				14'b01101100011111: oled_data = 16'b1111111111111111;
				14'b01101110011111: oled_data = 16'b1111111111111111;
				14'b01110000011111: oled_data = 16'b1111111111111111;
				14'b01110010011111: oled_data = 16'b1111111111111111;
				14'b01110100011111: oled_data = 16'b1111111111111111;
				14'b01110110011111: oled_data = 16'b1111111111111111;
				14'b01111000011111: oled_data = 16'b1111111111111111;
				14'b01111010011111: oled_data = 16'b1111111111111111;
				14'b01111100011111: oled_data = 16'b1111111111111111;
				14'b01111110011111: oled_data = 16'b1111111111111111;
				14'b10000000011111: oled_data = 16'b1111111111111111;
				14'b10000010011111: oled_data = 16'b1111111111111111;
				14'b10000100011111: oled_data = 16'b1111111111111111;
				14'b10000110011111: oled_data = 16'b1111111111111111;
				14'b10001000011111: oled_data = 16'b1111111111111111;
				14'b10001010011111: oled_data = 16'b1111111111111111;
				14'b10001100011111: oled_data = 16'b1111111111111111;
				14'b10001110011111: oled_data = 16'b1111111111111111;
				14'b10010000011111: oled_data = 16'b1111111111111111;
				14'b10010010011111: oled_data = 16'b1111111111111111;
				14'b10010100011111: oled_data = 16'b1111111111111111;
				14'b10010110011111: oled_data = 16'b1111111111111111;
				14'b10011000011111: oled_data = 16'b1111111111111111;
				14'b10011010011111: oled_data = 16'b1111111111111111;
				14'b10011100011111: oled_data = 16'b1111111111111111;
				14'b10011110011111: oled_data = 16'b1111111111111111;
				14'b10100000011111: oled_data = 16'b1111111111111111;
				14'b10100010011111: oled_data = 16'b1111111111111111;
				14'b10100100011111: oled_data = 16'b1111111111111111;
				14'b10100110011111: oled_data = 16'b1111111111111111;
				14'b10101000011111: oled_data = 16'b1111111111111111;
				14'b10101010011111: oled_data = 16'b1111111111111111;
				14'b10101100011111: oled_data = 16'b1111111111111111;
				14'b10101110011111: oled_data = 16'b1111111111111111;
				14'b10110000011111: oled_data = 16'b1111111111111111;
				14'b10110010011111: oled_data = 16'b1111111111111111;
				14'b10110100011111: oled_data = 16'b1111111111111111;
				14'b10110110011111: oled_data = 16'b1111111111111111;
				14'b10111000011111: oled_data = 16'b1111111111111111;
				14'b10111010011111: oled_data = 16'b1111111111111111;
				14'b10111100011111: oled_data = 16'b1111111111111111;
				14'b10111110011111: oled_data = 16'b1111111111111111;
				14'b00000000100000: oled_data = 16'b1111111111111111;
				14'b00000010100000: oled_data = 16'b1111111111111111;
				14'b00000100100000: oled_data = 16'b1111111111111111;
				14'b00000110100000: oled_data = 16'b1111111111111111;
				14'b00001000100000: oled_data = 16'b1111111111111111;
				14'b00001010100000: oled_data = 16'b1111111111111111;
				14'b00001100100000: oled_data = 16'b1111111111111111;
				14'b00001110100000: oled_data = 16'b1111111111111111;
				14'b00010000100000: oled_data = 16'b1111111111111111;
				14'b00010010100000: oled_data = 16'b1111111111111111;
				14'b00010100100000: oled_data = 16'b1111111111111111;
				14'b00010110100000: oled_data = 16'b1111111111111111;
				14'b00011000100000: oled_data = 16'b1111111111111111;
				14'b00011010100000: oled_data = 16'b1111111111111111;
				14'b00011100100000: oled_data = 16'b1111111111111111;
				14'b00011110100000: oled_data = 16'b1111111111111111;
				14'b00100000100000: oled_data = 16'b1111111111111111;
				14'b00100010100000: oled_data = 16'b1111111111111111;
				14'b00100100100000: oled_data = 16'b1111111111111111;
				14'b00100110100000: oled_data = 16'b1111111111111111;
				14'b00101000100000: oled_data = 16'b1111111111111111;
				14'b00101010100000: oled_data = 16'b1111111111111111;
				14'b00101100100000: oled_data = 16'b1111111111111111;
				14'b00101110100000: oled_data = 16'b1111111111111111;
				14'b00110000100000: oled_data = 16'b1111111111111111;
				14'b00110010100000: oled_data = 16'b1111111111111111;
				14'b00110100100000: oled_data = 16'b1111111111111111;
				14'b00110110100000: oled_data = 16'b1111111111111111;
				14'b00111000100000: oled_data = 16'b1111111111111111;
				14'b00111010100000: oled_data = 16'b1111111111111111;
				14'b00111100100000: oled_data = 16'b1111111111111111;
				14'b00111110100000: oled_data = 16'b1111111111111111;
				14'b01000000100000: oled_data = 16'b1111111111111111;
				14'b01000010100000: oled_data = 16'b1111111111111111;
				14'b01000100100000: oled_data = 16'b1111111111111111;
				14'b01000110100000: oled_data = 16'b1111111111111111;
				14'b01001000100000: oled_data = 16'b1111111111111111;
				14'b01001010100000: oled_data = 16'b1111111111111111;
				14'b01001100100000: oled_data = 16'b1111111111111111;
				14'b01001110100000: oled_data = 16'b1111111111111111;
				14'b01010000100000: oled_data = 16'b1111111111111111;
				14'b01010010100000: oled_data = 16'b1111111111111111;
				14'b01010100100000: oled_data = 16'b1111111111111111;
				14'b01010110100000: oled_data = 16'b1111111111111111;
				14'b01011000100000: oled_data = 16'b1111111111111111;
				14'b01011010100000: oled_data = 16'b1111111111111111;
				14'b01011100100000: oled_data = 16'b1111111111111111;
				14'b01011110100000: oled_data = 16'b1111111111111111;
				14'b01100000100000: oled_data = 16'b1111111111111111;
				14'b01100010100000: oled_data = 16'b1111111111111111;
				14'b01100100100000: oled_data = 16'b1111111111111111;
				14'b01100110100000: oled_data = 16'b1111111111111111;
				14'b01101000100000: oled_data = 16'b1111111111111111;
				14'b01101010100000: oled_data = 16'b1111111111111111;
				14'b01101100100000: oled_data = 16'b1111111111111111;
				14'b01101110100000: oled_data = 16'b1111111111111111;
				14'b01110000100000: oled_data = 16'b1111111111111111;
				14'b01110010100000: oled_data = 16'b1111111111111111;
				14'b01110100100000: oled_data = 16'b1111111111111111;
				14'b01110110100000: oled_data = 16'b1111111111111111;
				14'b01111000100000: oled_data = 16'b1111111111111111;
				14'b01111010100000: oled_data = 16'b1111111111111111;
				14'b01111100100000: oled_data = 16'b1111111111111111;
				14'b01111110100000: oled_data = 16'b1111111111111111;
				14'b10000000100000: oled_data = 16'b1111111111111111;
				14'b10000010100000: oled_data = 16'b1111111111111111;
				14'b10000100100000: oled_data = 16'b1111111111111111;
				14'b10000110100000: oled_data = 16'b1111111111111111;
				14'b10001000100000: oled_data = 16'b1111111111111111;
				14'b10001010100000: oled_data = 16'b1111111111111111;
				14'b10001100100000: oled_data = 16'b1111111111111111;
				14'b10001110100000: oled_data = 16'b1111111111111111;
				14'b10010000100000: oled_data = 16'b1111111111111111;
				14'b10010010100000: oled_data = 16'b1111111111111111;
				14'b10010100100000: oled_data = 16'b1111111111111111;
				14'b10010110100000: oled_data = 16'b1111111111111111;
				14'b10011000100000: oled_data = 16'b1111111111111111;
				14'b10011010100000: oled_data = 16'b1111111111111111;
				14'b10011100100000: oled_data = 16'b1111111111111111;
				14'b10011110100000: oled_data = 16'b1111111111111111;
				14'b10100000100000: oled_data = 16'b1111111111111111;
				14'b10100010100000: oled_data = 16'b1111111111111111;
				14'b10100100100000: oled_data = 16'b1111111111111111;
				14'b10100110100000: oled_data = 16'b1111111111111111;
				14'b10101000100000: oled_data = 16'b1111111111111111;
				14'b10101010100000: oled_data = 16'b1111111111111111;
				14'b10101100100000: oled_data = 16'b1111111111111111;
				14'b10101110100000: oled_data = 16'b1111111111111111;
				14'b10110000100000: oled_data = 16'b1111111111111111;
				14'b10110010100000: oled_data = 16'b1111111111111111;
				14'b10110100100000: oled_data = 16'b1111111111111111;
				14'b10110110100000: oled_data = 16'b1111111111111111;
				14'b10111000100000: oled_data = 16'b1111111111111111;
				14'b10111010100000: oled_data = 16'b1111111111111111;
				14'b10111100100000: oled_data = 16'b1111111111111111;
				14'b10111110100000: oled_data = 16'b1111111111111111;
				14'b00000000100001: oled_data = 16'b1111111111111111;
				14'b00000010100001: oled_data = 16'b1111111111111111;
				14'b00000100100001: oled_data = 16'b1111111111111111;
				14'b00000110100001: oled_data = 16'b1111111111111111;
				14'b00001000100001: oled_data = 16'b1111111111111111;
				14'b00001010100001: oled_data = 16'b1111111111111111;
				14'b00001100100001: oled_data = 16'b1111111111111111;
				14'b00001110100001: oled_data = 16'b1111111111111111;
				14'b00010000100001: oled_data = 16'b1111111111111111;
				14'b00010010100001: oled_data = 16'b1111111111111111;
				14'b00010100100001: oled_data = 16'b1111111111111111;
				14'b00010110100001: oled_data = 16'b1111111111111111;
				14'b00011000100001: oled_data = 16'b1111111111111111;
				14'b00011010100001: oled_data = 16'b1111111111111111;
				14'b00011100100001: oled_data = 16'b1111111111111111;
				14'b00011110100001: oled_data = 16'b1111111111111111;
				14'b00100000100001: oled_data = 16'b1111111111111111;
				14'b00100010100001: oled_data = 16'b1111111111111111;
				14'b00100100100001: oled_data = 16'b1111111111111111;
				14'b00100110100001: oled_data = 16'b1111111111111111;
				14'b00101000100001: oled_data = 16'b1111111111111111;
				14'b00101010100001: oled_data = 16'b1111111111111111;
				14'b00101100100001: oled_data = 16'b1111111111111111;
				14'b00101110100001: oled_data = 16'b1111111111111111;
				14'b00110000100001: oled_data = 16'b1111111111111111;
				14'b00110010100001: oled_data = 16'b1111111111111111;
				14'b00110100100001: oled_data = 16'b1111111111111111;
				14'b00110110100001: oled_data = 16'b1111111111111111;
				14'b00111000100001: oled_data = 16'b1111111111111111;
				14'b00111010100001: oled_data = 16'b1111111111111111;
				14'b00111100100001: oled_data = 16'b1111111111111111;
				14'b00111110100001: oled_data = 16'b1111111111111111;
				14'b01000000100001: oled_data = 16'b1111111111111111;
				14'b01000010100001: oled_data = 16'b1111111111111111;
				14'b01000100100001: oled_data = 16'b1111111111111111;
				14'b01000110100001: oled_data = 16'b1111111111111111;
				14'b01001000100001: oled_data = 16'b1111111111111111;
				14'b01001010100001: oled_data = 16'b1111111111111111;
				14'b01001100100001: oled_data = 16'b1111111111111111;
				14'b01001110100001: oled_data = 16'b1111111111111111;
				14'b01010000100001: oled_data = 16'b1111111111111111;
				14'b01010010100001: oled_data = 16'b1111111111111111;
				14'b01010100100001: oled_data = 16'b1111111111111111;
				14'b01010110100001: oled_data = 16'b1111111111111111;
				14'b01011000100001: oled_data = 16'b1111111111111111;
				14'b01011010100001: oled_data = 16'b1111111111111111;
				14'b01011100100001: oled_data = 16'b1111111111111111;
				14'b01011110100001: oled_data = 16'b1111111111111111;
				14'b01100000100001: oled_data = 16'b1111111111111111;
				14'b01100010100001: oled_data = 16'b1111111111111111;
				14'b01100100100001: oled_data = 16'b1111111111111111;
				14'b01100110100001: oled_data = 16'b1111111111111111;
				14'b01101000100001: oled_data = 16'b1111111111111111;
				14'b01101010100001: oled_data = 16'b1111111111111111;
				14'b01101100100001: oled_data = 16'b1111111111111111;
				14'b01101110100001: oled_data = 16'b1111111111111111;
				14'b01110000100001: oled_data = 16'b1111111111111111;
				14'b01110010100001: oled_data = 16'b1111111111111111;
				14'b01110100100001: oled_data = 16'b1111111111111111;
				14'b01110110100001: oled_data = 16'b1111111111111111;
				14'b01111000100001: oled_data = 16'b1111111111111111;
				14'b01111010100001: oled_data = 16'b1111111111111111;
				14'b01111100100001: oled_data = 16'b1111111111111111;
				14'b01111110100001: oled_data = 16'b1111111111111111;
				14'b10000000100001: oled_data = 16'b1111111111111111;
				14'b10000010100001: oled_data = 16'b1111111111111111;
				14'b10000100100001: oled_data = 16'b1111111111111111;
				14'b10000110100001: oled_data = 16'b1111111111111111;
				14'b10001000100001: oled_data = 16'b1111111111111111;
				14'b10001010100001: oled_data = 16'b1111111111111111;
				14'b10001100100001: oled_data = 16'b1111111111111111;
				14'b10001110100001: oled_data = 16'b1111111111111111;
				14'b10010000100001: oled_data = 16'b1111111111111111;
				14'b10010010100001: oled_data = 16'b1111111111111111;
				14'b10010100100001: oled_data = 16'b1111111111111111;
				14'b10010110100001: oled_data = 16'b1111111111111111;
				14'b10011000100001: oled_data = 16'b1111111111111111;
				14'b10011010100001: oled_data = 16'b1111111111111111;
				14'b10011100100001: oled_data = 16'b1111111111111111;
				14'b10011110100001: oled_data = 16'b1111111111111111;
				14'b10100000100001: oled_data = 16'b1111111111111111;
				14'b10100010100001: oled_data = 16'b1111111111111111;
				14'b10100100100001: oled_data = 16'b1111111111111111;
				14'b10100110100001: oled_data = 16'b1111111111111111;
				14'b10101000100001: oled_data = 16'b1111111111111111;
				14'b10101010100001: oled_data = 16'b1111111111111111;
				14'b10101100100001: oled_data = 16'b1111111111111111;
				14'b10101110100001: oled_data = 16'b1111111111111111;
				14'b10110000100001: oled_data = 16'b1111111111111111;
				14'b10110010100001: oled_data = 16'b1111111111111111;
				14'b10110100100001: oled_data = 16'b1111111111111111;
				14'b10110110100001: oled_data = 16'b1111111111111111;
				14'b10111000100001: oled_data = 16'b1111111111111111;
				14'b10111010100001: oled_data = 16'b1111111111111111;
				14'b10111100100001: oled_data = 16'b1111111111111111;
				14'b10111110100001: oled_data = 16'b1111111111111111;
				14'b00000000100010: oled_data = 16'b1111111111111111;
				14'b00000010100010: oled_data = 16'b1111111111111111;
				14'b00000100100010: oled_data = 16'b1111111111111111;
				14'b00000110100010: oled_data = 16'b1111111111111111;
				14'b00001000100010: oled_data = 16'b1111111111111111;
				14'b00001010100010: oled_data = 16'b1111111111111111;
				14'b00001100100010: oled_data = 16'b1111111111111111;
				14'b00001110100010: oled_data = 16'b1111111111111111;
				14'b00010000100010: oled_data = 16'b1111111111111111;
				14'b00010010100010: oled_data = 16'b1111111111111111;
				14'b00010100100010: oled_data = 16'b1111111111111111;
				14'b00010110100010: oled_data = 16'b1111111111111111;
				14'b00011000100010: oled_data = 16'b1111111111111111;
				14'b00011010100010: oled_data = 16'b1111111111111111;
				14'b00011100100010: oled_data = 16'b1111111111111111;
				14'b00011110100010: oled_data = 16'b1111111111111111;
				14'b00100000100010: oled_data = 16'b1111111111111111;
				14'b00100010100010: oled_data = 16'b1111111111111111;
				14'b00100100100010: oled_data = 16'b1111111111111111;
				14'b00100110100010: oled_data = 16'b1111111111111111;
				14'b00101000100010: oled_data = 16'b1111111111111111;
				14'b00101010100010: oled_data = 16'b1111111111111111;
				14'b00101100100010: oled_data = 16'b1111111111111111;
				14'b00101110100010: oled_data = 16'b1111111111111111;
				14'b00110000100010: oled_data = 16'b1111111111111111;
				14'b00110010100010: oled_data = 16'b1111111111111111;
				14'b00110100100010: oled_data = 16'b1111111111111111;
				14'b00110110100010: oled_data = 16'b1111111111111111;
				14'b00111000100010: oled_data = 16'b1111111111111111;
				14'b00111010100010: oled_data = 16'b1111111111111111;
				14'b00111100100010: oled_data = 16'b1111111111111111;
				14'b00111110100010: oled_data = 16'b1111111111111111;
				14'b01000000100010: oled_data = 16'b1111111111111111;
				14'b01000010100010: oled_data = 16'b1111111111111111;
				14'b01000100100010: oled_data = 16'b1111111111111111;
				14'b01000110100010: oled_data = 16'b1111111111111111;
				14'b01001000100010: oled_data = 16'b1111111111111111;
				14'b01001010100010: oled_data = 16'b1111111111111111;
				14'b01001100100010: oled_data = 16'b1111111111111111;
				14'b01001110100010: oled_data = 16'b1111111111111111;
				14'b01010000100010: oled_data = 16'b1111111111111111;
				14'b01010010100010: oled_data = 16'b1111111111111111;
				14'b01010100100010: oled_data = 16'b1111111111111111;
				14'b01010110100010: oled_data = 16'b1111111111111111;
				14'b01011000100010: oled_data = 16'b1111111111111111;
				14'b01011010100010: oled_data = 16'b1111111111111111;
				14'b01011100100010: oled_data = 16'b1111111111111111;
				14'b01011110100010: oled_data = 16'b1111111111111111;
				14'b01100000100010: oled_data = 16'b1111111111111111;
				14'b01100010100010: oled_data = 16'b1111111111111111;
				14'b01100100100010: oled_data = 16'b1111111111111111;
				14'b01100110100010: oled_data = 16'b1111111111111111;
				14'b01101000100010: oled_data = 16'b1111111111111111;
				14'b01101010100010: oled_data = 16'b1111111111111111;
				14'b01101100100010: oled_data = 16'b1111111111111111;
				14'b01101110100010: oled_data = 16'b1111111111111111;
				14'b01110000100010: oled_data = 16'b1111111111111111;
				14'b01110010100010: oled_data = 16'b1111111111111111;
				14'b01110100100010: oled_data = 16'b1111111111111111;
				14'b01110110100010: oled_data = 16'b1111111111111111;
				14'b01111000100010: oled_data = 16'b1111111111111111;
				14'b01111010100010: oled_data = 16'b1111111111111111;
				14'b01111100100010: oled_data = 16'b1111111111111111;
				14'b01111110100010: oled_data = 16'b1111111111111111;
				14'b10000000100010: oled_data = 16'b1111111111111111;
				14'b10000010100010: oled_data = 16'b1111111111111111;
				14'b10000100100010: oled_data = 16'b1111111111111111;
				14'b10000110100010: oled_data = 16'b1111111111111111;
				14'b10001000100010: oled_data = 16'b1111111111111111;
				14'b10001010100010: oled_data = 16'b1111111111111111;
				14'b10001100100010: oled_data = 16'b1111111111111111;
				14'b10001110100010: oled_data = 16'b1111111111111111;
				14'b10010000100010: oled_data = 16'b1111111111111111;
				14'b10010010100010: oled_data = 16'b1111111111111111;
				14'b10010100100010: oled_data = 16'b1111111111111111;
				14'b10010110100010: oled_data = 16'b1111111111111111;
				14'b10011000100010: oled_data = 16'b1111111111111111;
				14'b10011010100010: oled_data = 16'b1111111111111111;
				14'b10011100100010: oled_data = 16'b1111111111111111;
				14'b10011110100010: oled_data = 16'b1111111111111111;
				14'b10100000100010: oled_data = 16'b1111111111111111;
				14'b10100010100010: oled_data = 16'b1111111111111111;
				14'b10100100100010: oled_data = 16'b1111111111111111;
				14'b10100110100010: oled_data = 16'b1111111111111111;
				14'b10101000100010: oled_data = 16'b1111111111111111;
				14'b10101010100010: oled_data = 16'b1111111111111111;
				14'b10101100100010: oled_data = 16'b1111111111111111;
				14'b10101110100010: oled_data = 16'b1111111111111111;
				14'b10110000100010: oled_data = 16'b1111111111111111;
				14'b10110010100010: oled_data = 16'b1111111111111111;
				14'b10110100100010: oled_data = 16'b1111111111111111;
				14'b10110110100010: oled_data = 16'b1111111111111111;
				14'b10111000100010: oled_data = 16'b1111111111111111;
				14'b10111010100010: oled_data = 16'b1111111111111111;
				14'b10111100100010: oled_data = 16'b1111111111111111;
				14'b10111110100010: oled_data = 16'b1111111111111111;
				14'b00000000100011: oled_data = 16'b1111111111111111;
				14'b00000010100011: oled_data = 16'b1111111111111111;
				14'b00000100100011: oled_data = 16'b1111111111111111;
				14'b00000110100011: oled_data = 16'b1111111111111111;
				14'b00001000100011: oled_data = 16'b1111111111111111;
				14'b00001010100011: oled_data = 16'b1111111111111111;
				14'b00001100100011: oled_data = 16'b1111111111111111;
				14'b00001110100011: oled_data = 16'b1111111111111111;
				14'b00010000100011: oled_data = 16'b1111111111111111;
				14'b00010010100011: oled_data = 16'b1111111111111111;
				14'b00010100100011: oled_data = 16'b1111111111111111;
				14'b00010110100011: oled_data = 16'b1111111111111111;
				14'b00011000100011: oled_data = 16'b1111111111111111;
				14'b00011010100011: oled_data = 16'b1111111111111111;
				14'b00011100100011: oled_data = 16'b1111111111111111;
				14'b00011110100011: oled_data = 16'b1111111111111111;
				14'b00100000100011: oled_data = 16'b1111111111111111;
				14'b00100010100011: oled_data = 16'b1111111111111111;
				14'b00100100100011: oled_data = 16'b1111111111111111;
				14'b00100110100011: oled_data = 16'b1111111111111111;
				14'b00101000100011: oled_data = 16'b1111111111111111;
				14'b00101010100011: oled_data = 16'b1111111111111111;
				14'b00101100100011: oled_data = 16'b1111111111111111;
				14'b00101110100011: oled_data = 16'b1111111111111111;
				14'b00110000100011: oled_data = 16'b1111111111111111;
				14'b00110010100011: oled_data = 16'b1111111111111111;
				14'b00110100100011: oled_data = 16'b1111111111111111;
				14'b00110110100011: oled_data = 16'b1111111111111111;
				14'b00111000100011: oled_data = 16'b1111111111111111;
				14'b00111010100011: oled_data = 16'b1111111111111111;
				14'b00111100100011: oled_data = 16'b1111111111111111;
				14'b00111110100011: oled_data = 16'b1111111111111111;
				14'b01000000100011: oled_data = 16'b1111111111111111;
				14'b01000010100011: oled_data = 16'b1111111111111111;
				14'b01000100100011: oled_data = 16'b1111111111111111;
				14'b01000110100011: oled_data = 16'b1111111111111111;
				14'b01001000100011: oled_data = 16'b1111111111111111;
				14'b01001010100011: oled_data = 16'b1111111111111111;
				14'b01001100100011: oled_data = 16'b1111111111111111;
				14'b01001110100011: oled_data = 16'b1111111111111111;
				14'b01010000100011: oled_data = 16'b1111111111111111;
				14'b01010010100011: oled_data = 16'b1111111111111111;
				14'b01010100100011: oled_data = 16'b1111111111111111;
				14'b01010110100011: oled_data = 16'b1111111111111111;
				14'b01011000100011: oled_data = 16'b1111111111111111;
				14'b01011010100011: oled_data = 16'b1111111111111111;
				14'b01011100100011: oled_data = 16'b1111111111111111;
				14'b01011110100011: oled_data = 16'b1111111111111111;
				14'b01100000100011: oled_data = 16'b1111111111111111;
				14'b01100010100011: oled_data = 16'b1111111111111111;
				14'b01100100100011: oled_data = 16'b1111111111111111;
				14'b01100110100011: oled_data = 16'b1111111111111111;
				14'b01101000100011: oled_data = 16'b1111111111111111;
				14'b01101010100011: oled_data = 16'b1111111111111111;
				14'b01101100100011: oled_data = 16'b1111111111111111;
				14'b01101110100011: oled_data = 16'b1111111111111111;
				14'b01110000100011: oled_data = 16'b1111111111111111;
				14'b01110010100011: oled_data = 16'b1111111111111111;
				14'b01110100100011: oled_data = 16'b1111111111111111;
				14'b01110110100011: oled_data = 16'b1111111111111111;
				14'b01111000100011: oled_data = 16'b1111111111111111;
				14'b01111010100011: oled_data = 16'b1111111111111111;
				14'b01111100100011: oled_data = 16'b1111111111111111;
				14'b01111110100011: oled_data = 16'b1111111111111111;
				14'b10000000100011: oled_data = 16'b1111111111111111;
				14'b10000010100011: oled_data = 16'b1111111111111111;
				14'b10000100100011: oled_data = 16'b1111111111111111;
				14'b10000110100011: oled_data = 16'b1111111111111111;
				14'b10001000100011: oled_data = 16'b1111111111111111;
				14'b10001010100011: oled_data = 16'b1111111111111111;
				14'b10001100100011: oled_data = 16'b1111111111111111;
				14'b10001110100011: oled_data = 16'b1111111111111111;
				14'b10010000100011: oled_data = 16'b1111111111111111;
				14'b10010010100011: oled_data = 16'b1111111111111111;
				14'b10010100100011: oled_data = 16'b1111111111111111;
				14'b10010110100011: oled_data = 16'b1111111111111111;
				14'b10011000100011: oled_data = 16'b1111111111111111;
				14'b10011010100011: oled_data = 16'b1111111111111111;
				14'b10011100100011: oled_data = 16'b1111111111111111;
				14'b10011110100011: oled_data = 16'b1111111111111111;
				14'b10100000100011: oled_data = 16'b1111111111111111;
				14'b10100010100011: oled_data = 16'b1111111111111111;
				14'b10100100100011: oled_data = 16'b1111111111111111;
				14'b10100110100011: oled_data = 16'b1111111111111111;
				14'b10101000100011: oled_data = 16'b1111111111111111;
				14'b10101010100011: oled_data = 16'b1111111111111111;
				14'b10101100100011: oled_data = 16'b1111111111111111;
				14'b10101110100011: oled_data = 16'b1111111111111111;
				14'b10110000100011: oled_data = 16'b1111111111111111;
				14'b10110010100011: oled_data = 16'b1111111111111111;
				14'b10110100100011: oled_data = 16'b1111111111111111;
				14'b10110110100011: oled_data = 16'b1111111111111111;
				14'b10111000100011: oled_data = 16'b1111111111111111;
				14'b10111010100011: oled_data = 16'b1111111111111111;
				14'b10111100100011: oled_data = 16'b1111111111111111;
				14'b10111110100011: oled_data = 16'b1111111111111111;
				14'b00000000100100: oled_data = 16'b1111111111111111;
				14'b00000010100100: oled_data = 16'b1111111111111111;
				14'b00000100100100: oled_data = 16'b1111111111111111;
				14'b00000110100100: oled_data = 16'b1111111111111111;
				14'b00001000100100: oled_data = 16'b1111111111111111;
				14'b00001010100100: oled_data = 16'b1111111111111111;
				14'b00001100100100: oled_data = 16'b1111111111111111;
				14'b00001110100100: oled_data = 16'b1111111111111111;
				14'b00010000100100: oled_data = 16'b1111111111111111;
				14'b00010010100100: oled_data = 16'b1111111111111111;
				14'b00010100100100: oled_data = 16'b1111111111111111;
				14'b00010110100100: oled_data = 16'b1111111111111111;
				14'b00011000100100: oled_data = 16'b1111111111111111;
				14'b00011010100100: oled_data = 16'b1111111111111111;
				14'b00011100100100: oled_data = 16'b1111111111111111;
				14'b00011110100100: oled_data = 16'b1111111111111111;
				14'b00100000100100: oled_data = 16'b1111111111111111;
				14'b00100010100100: oled_data = 16'b1111111111111111;
				14'b00100100100100: oled_data = 16'b1111111111111111;
				14'b00100110100100: oled_data = 16'b1111111111111111;
				14'b00101000100100: oled_data = 16'b1111111111111111;
				14'b00101010100100: oled_data = 16'b1111111111111111;
				14'b00101100100100: oled_data = 16'b1111111111111111;
				14'b00101110100100: oled_data = 16'b1111111111111111;
				14'b00110000100100: oled_data = 16'b1111111111111111;
				14'b00110010100100: oled_data = 16'b1111111111111111;
				14'b00110100100100: oled_data = 16'b1111111111111111;
				14'b00110110100100: oled_data = 16'b1111111111111111;
				14'b00111000100100: oled_data = 16'b1111111111111111;
				14'b00111010100100: oled_data = 16'b1111111111111111;
				14'b00111100100100: oled_data = 16'b1111111111111111;
				14'b00111110100100: oled_data = 16'b1111111111111111;
				14'b01000000100100: oled_data = 16'b1111111111111111;
				14'b01000010100100: oled_data = 16'b1111111111111111;
				14'b01000100100100: oled_data = 16'b1111111111111111;
				14'b01000110100100: oled_data = 16'b1111111111111111;
				14'b01001000100100: oled_data = 16'b1111111111111111;
				14'b01001010100100: oled_data = 16'b1111111111111111;
				14'b01001100100100: oled_data = 16'b1111111111111111;
				14'b01001110100100: oled_data = 16'b1111111111111111;
				14'b01010000100100: oled_data = 16'b1111111111111111;
				14'b01010010100100: oled_data = 16'b1111111111111111;
				14'b01010100100100: oled_data = 16'b1111111111111111;
				14'b01010110100100: oled_data = 16'b1111111111111111;
				14'b01011000100100: oled_data = 16'b1111111111111111;
				14'b01011010100100: oled_data = 16'b1111111111111111;
				14'b01011100100100: oled_data = 16'b1111111111111111;
				14'b01011110100100: oled_data = 16'b1111111111111111;
				14'b01100000100100: oled_data = 16'b1111111111111111;
				14'b01100010100100: oled_data = 16'b1111111111111111;
				14'b01100100100100: oled_data = 16'b1111111111111111;
				14'b01100110100100: oled_data = 16'b1111111111111111;
				14'b01101000100100: oled_data = 16'b1111111111111111;
				14'b01101010100100: oled_data = 16'b1111111111111111;
				14'b01101100100100: oled_data = 16'b1111111111111111;
				14'b01101110100100: oled_data = 16'b1111111111111111;
				14'b01110000100100: oled_data = 16'b1111111111111111;
				14'b01110010100100: oled_data = 16'b1111111111111111;
				14'b01110100100100: oled_data = 16'b1111111111111111;
				14'b01110110100100: oled_data = 16'b1111111111111111;
				14'b01111000100100: oled_data = 16'b1111111111111111;
				14'b01111010100100: oled_data = 16'b1111111111111111;
				14'b01111100100100: oled_data = 16'b1111111111111111;
				14'b01111110100100: oled_data = 16'b1111111111111111;
				14'b10000000100100: oled_data = 16'b1111111111111111;
				14'b10000010100100: oled_data = 16'b1111111111111111;
				14'b10000100100100: oled_data = 16'b1111111111111111;
				14'b10000110100100: oled_data = 16'b1111111111111111;
				14'b10001000100100: oled_data = 16'b1111111111111111;
				14'b10001010100100: oled_data = 16'b1111111111111111;
				14'b10001100100100: oled_data = 16'b1111111111111111;
				14'b10001110100100: oled_data = 16'b1111111111111111;
				14'b10010000100100: oled_data = 16'b1111111111111111;
				14'b10010010100100: oled_data = 16'b1111111111111111;
				14'b10010100100100: oled_data = 16'b1111111111111111;
				14'b10010110100100: oled_data = 16'b1111111111111111;
				14'b10011000100100: oled_data = 16'b1111111111111111;
				14'b10011010100100: oled_data = 16'b1111111111111111;
				14'b10011100100100: oled_data = 16'b1111111111111111;
				14'b10011110100100: oled_data = 16'b1111111111111111;
				14'b10100000100100: oled_data = 16'b1111111111111111;
				14'b10100010100100: oled_data = 16'b1111111111111111;
				14'b10100100100100: oled_data = 16'b1111111111111111;
				14'b10100110100100: oled_data = 16'b1111111111111111;
				14'b10101000100100: oled_data = 16'b1111111111111111;
				14'b10101010100100: oled_data = 16'b1111111111111111;
				14'b10101100100100: oled_data = 16'b1111111111111111;
				14'b10101110100100: oled_data = 16'b1111111111111111;
				14'b10110000100100: oled_data = 16'b1111111111111111;
				14'b10110010100100: oled_data = 16'b1111111111111111;
				14'b10110100100100: oled_data = 16'b1111111111111111;
				14'b10110110100100: oled_data = 16'b1111111111111111;
				14'b10111000100100: oled_data = 16'b1111111111111111;
				14'b10111010100100: oled_data = 16'b1111111111111111;
				14'b10111100100100: oled_data = 16'b1111111111111111;
				14'b10111110100100: oled_data = 16'b1111111111111111;
				14'b00000000100101: oled_data = 16'b1111111111111111;
				14'b00000010100101: oled_data = 16'b1111111111111111;
				14'b00000100100101: oled_data = 16'b1111111111111111;
				14'b00000110100101: oled_data = 16'b1111111111111111;
				14'b00001000100101: oled_data = 16'b1111111111111111;
				14'b00001010100101: oled_data = 16'b1111111111111111;
				14'b00001100100101: oled_data = 16'b1111111111111111;
				14'b00001110100101: oled_data = 16'b1111111111111111;
				14'b00010000100101: oled_data = 16'b1111111111111111;
				14'b00010010100101: oled_data = 16'b1111111111111111;
				14'b00010100100101: oled_data = 16'b1111111111111111;
				14'b00010110100101: oled_data = 16'b1111111111111111;
				14'b00011000100101: oled_data = 16'b1111111111111111;
				14'b00011010100101: oled_data = 16'b1111111111111111;
				14'b00011100100101: oled_data = 16'b1111111111111111;
				14'b00011110100101: oled_data = 16'b1111111111111111;
				14'b00100000100101: oled_data = 16'b1111111111111111;
				14'b00100010100101: oled_data = 16'b1111111111111111;
				14'b00100100100101: oled_data = 16'b1111111111111111;
				14'b00100110100101: oled_data = 16'b1111111111111111;
				14'b00101000100101: oled_data = 16'b1111111111111111;
				14'b00101010100101: oled_data = 16'b1111111111111111;
				14'b00101100100101: oled_data = 16'b1111111111111111;
				14'b00101110100101: oled_data = 16'b1111111111111111;
				14'b00110000100101: oled_data = 16'b1111111111111111;
				14'b00110010100101: oled_data = 16'b1111111111111111;
				14'b00110100100101: oled_data = 16'b1111111111111111;
				14'b00110110100101: oled_data = 16'b1111111111111111;
				14'b00111000100101: oled_data = 16'b1111111111111111;
				14'b00111010100101: oled_data = 16'b1111111111111111;
				14'b00111100100101: oled_data = 16'b1111111111111111;
				14'b00111110100101: oled_data = 16'b1111111111111111;
				14'b01000000100101: oled_data = 16'b1111111111111111;
				14'b01000010100101: oled_data = 16'b1111111111111111;
				14'b01000100100101: oled_data = 16'b1111111111111111;
				14'b01000110100101: oled_data = 16'b1111111111111111;
				14'b01001000100101: oled_data = 16'b1111111111111111;
				14'b01001010100101: oled_data = 16'b1111111111111111;
				14'b01001100100101: oled_data = 16'b1111111111111111;
				14'b01001110100101: oled_data = 16'b1111111111111111;
				14'b01010000100101: oled_data = 16'b1111111111111111;
				14'b01010010100101: oled_data = 16'b1111111111111111;
				14'b01010100100101: oled_data = 16'b1111111111111111;
				14'b01010110100101: oled_data = 16'b1111111111111111;
				14'b01011000100101: oled_data = 16'b1111111111111111;
				14'b01011010100101: oled_data = 16'b1111111111111111;
				14'b01011100100101: oled_data = 16'b1111111111111111;
				14'b01011110100101: oled_data = 16'b1111111111111111;
				14'b01100000100101: oled_data = 16'b1111111111111111;
				14'b01100010100101: oled_data = 16'b1111111111111111;
				14'b01100100100101: oled_data = 16'b1111111111111111;
				14'b01100110100101: oled_data = 16'b1111111111111111;
				14'b01101000100101: oled_data = 16'b1111111111111111;
				14'b01101010100101: oled_data = 16'b1111111111111111;
				14'b01101100100101: oled_data = 16'b1111111111111111;
				14'b01101110100101: oled_data = 16'b1111111111111111;
				14'b01110000100101: oled_data = 16'b1111111111111111;
				14'b01110010100101: oled_data = 16'b1111111111111111;
				14'b01110100100101: oled_data = 16'b1111111111111111;
				14'b01110110100101: oled_data = 16'b1111111111111111;
				14'b01111000100101: oled_data = 16'b1111111111111111;
				14'b01111010100101: oled_data = 16'b1111111111111111;
				14'b01111100100101: oled_data = 16'b1111111111111111;
				14'b01111110100101: oled_data = 16'b1111111111111111;
				14'b10000000100101: oled_data = 16'b1111111111111111;
				14'b10000010100101: oled_data = 16'b1111111111111111;
				14'b10000100100101: oled_data = 16'b1111111111111111;
				14'b10000110100101: oled_data = 16'b1111111111111111;
				14'b10001000100101: oled_data = 16'b1111111111111111;
				14'b10001010100101: oled_data = 16'b1111111111111111;
				14'b10001100100101: oled_data = 16'b1111111111111111;
				14'b10001110100101: oled_data = 16'b1111111111111111;
				14'b10010000100101: oled_data = 16'b1111111111111111;
				14'b10010010100101: oled_data = 16'b1111111111111111;
				14'b10010100100101: oled_data = 16'b1111111111111111;
				14'b10010110100101: oled_data = 16'b1111111111111111;
				14'b10011000100101: oled_data = 16'b1111111111111111;
				14'b10011010100101: oled_data = 16'b1111111111111111;
				14'b10011100100101: oled_data = 16'b1111111111111111;
				14'b10011110100101: oled_data = 16'b1111111111111111;
				14'b10100000100101: oled_data = 16'b1111111111111111;
				14'b10100010100101: oled_data = 16'b1111111111111111;
				14'b10100100100101: oled_data = 16'b1111111111111111;
				14'b10100110100101: oled_data = 16'b1111111111111111;
				14'b10101000100101: oled_data = 16'b1111111111111111;
				14'b10101010100101: oled_data = 16'b1111111111111111;
				14'b10101100100101: oled_data = 16'b1111111111111111;
				14'b10101110100101: oled_data = 16'b1111111111111111;
				14'b10110000100101: oled_data = 16'b1111111111111111;
				14'b10110010100101: oled_data = 16'b1111111111111111;
				14'b10110100100101: oled_data = 16'b1111111111111111;
				14'b10110110100101: oled_data = 16'b1111111111111111;
				14'b10111000100101: oled_data = 16'b1111111111111111;
				14'b10111010100101: oled_data = 16'b1111111111111111;
				14'b10111100100101: oled_data = 16'b1111111111111111;
				14'b10111110100101: oled_data = 16'b1111111111111111;
				14'b00000000100110: oled_data = 16'b1111111111111111;
				14'b00000010100110: oled_data = 16'b1111111111111111;
				14'b00000100100110: oled_data = 16'b1111111111111111;
				14'b00000110100110: oled_data = 16'b1111111111111111;
				14'b00001000100110: oled_data = 16'b1111111111111111;
				14'b00001010100110: oled_data = 16'b1111111111111111;
				14'b00001100100110: oled_data = 16'b1111111111111111;
				14'b00001110100110: oled_data = 16'b1111111111111111;
				14'b00010000100110: oled_data = 16'b1111111111111111;
				14'b00010010100110: oled_data = 16'b1111111111111111;
				14'b00010100100110: oled_data = 16'b1111111111111111;
				14'b00010110100110: oled_data = 16'b1111111111111111;
				14'b00011000100110: oled_data = 16'b1111111111111111;
				14'b00011010100110: oled_data = 16'b1111111111111111;
				14'b00011100100110: oled_data = 16'b1111111111111111;
				14'b00011110100110: oled_data = 16'b1111111111111111;
				14'b00100000100110: oled_data = 16'b1111111111111111;
				14'b00100010100110: oled_data = 16'b1111111111111111;
				14'b00100100100110: oled_data = 16'b1111111111111111;
				14'b00100110100110: oled_data = 16'b1111111111111111;
				14'b00101000100110: oled_data = 16'b1111111111111111;
				14'b00101010100110: oled_data = 16'b1111111111111111;
				14'b00101100100110: oled_data = 16'b1111111111111111;
				14'b00101110100110: oled_data = 16'b1111111111111111;
				14'b00110000100110: oled_data = 16'b1111111111111111;
				14'b00110010100110: oled_data = 16'b1111111111111111;
				14'b00110100100110: oled_data = 16'b1111111111111111;
				14'b00110110100110: oled_data = 16'b1111111111111111;
				14'b00111000100110: oled_data = 16'b1111111111111111;
				14'b00111010100110: oled_data = 16'b1111111111111111;
				14'b00111100100110: oled_data = 16'b1111111111111111;
				14'b00111110100110: oled_data = 16'b1111111111111111;
				14'b01000000100110: oled_data = 16'b1111111111111111;
				14'b01000010100110: oled_data = 16'b1111111111111111;
				14'b01000100100110: oled_data = 16'b1111111111111111;
				14'b01000110100110: oled_data = 16'b1111111111111111;
				14'b01001000100110: oled_data = 16'b1111111111111111;
				14'b01001010100110: oled_data = 16'b1111111111111111;
				14'b01001100100110: oled_data = 16'b1111111111111111;
				14'b01001110100110: oled_data = 16'b1111111111111111;
				14'b01010000100110: oled_data = 16'b1111111111111111;
				14'b01010010100110: oled_data = 16'b1111111111111111;
				14'b01010100100110: oled_data = 16'b1111111111111111;
				14'b01010110100110: oled_data = 16'b1111111111111111;
				14'b01011000100110: oled_data = 16'b1111111111111111;
				14'b01011010100110: oled_data = 16'b1111111111111111;
				14'b01011100100110: oled_data = 16'b1111111111111111;
				14'b01011110100110: oled_data = 16'b1111111111111111;
				14'b01100000100110: oled_data = 16'b1111111111111111;
				14'b01100010100110: oled_data = 16'b1111111111111111;
				14'b01100100100110: oled_data = 16'b1111111111111111;
				14'b01100110100110: oled_data = 16'b1111111111111111;
				14'b01101000100110: oled_data = 16'b1111111111111111;
				14'b01101010100110: oled_data = 16'b1111111111111111;
				14'b01101100100110: oled_data = 16'b1111111111111111;
				14'b01101110100110: oled_data = 16'b1111111111111111;
				14'b01110000100110: oled_data = 16'b1111111111111111;
				14'b01110010100110: oled_data = 16'b1111111111111111;
				14'b01110100100110: oled_data = 16'b1111111111111111;
				14'b01110110100110: oled_data = 16'b1111111111111111;
				14'b01111000100110: oled_data = 16'b1111111111111111;
				14'b01111010100110: oled_data = 16'b1111111111111111;
				14'b01111100100110: oled_data = 16'b1111111111111111;
				14'b01111110100110: oled_data = 16'b1111111111111111;
				14'b10000000100110: oled_data = 16'b1111111111111111;
				14'b10000010100110: oled_data = 16'b1111111111111111;
				14'b10000100100110: oled_data = 16'b1111111111111111;
				14'b10000110100110: oled_data = 16'b1111111111111111;
				14'b10001000100110: oled_data = 16'b1111111111111111;
				14'b10001010100110: oled_data = 16'b1111111111111111;
				14'b10001100100110: oled_data = 16'b1111111111111111;
				14'b10001110100110: oled_data = 16'b1111111111111111;
				14'b10010000100110: oled_data = 16'b1111111111111111;
				14'b10010010100110: oled_data = 16'b1111111111111111;
				14'b10010100100110: oled_data = 16'b1111111111111111;
				14'b10010110100110: oled_data = 16'b1111111111111111;
				14'b10011000100110: oled_data = 16'b1111111111111111;
				14'b10011010100110: oled_data = 16'b1111111111111111;
				14'b10011100100110: oled_data = 16'b1111111111111111;
				14'b10011110100110: oled_data = 16'b1111111111111111;
				14'b10100000100110: oled_data = 16'b1111111111111111;
				14'b10100010100110: oled_data = 16'b1111111111111111;
				14'b10100100100110: oled_data = 16'b1111111111111111;
				14'b10100110100110: oled_data = 16'b1111111111111111;
				14'b10101000100110: oled_data = 16'b1111111111111111;
				14'b10101010100110: oled_data = 16'b1111111111111111;
				14'b10101100100110: oled_data = 16'b1111111111111111;
				14'b10101110100110: oled_data = 16'b1111111111111111;
				14'b10110000100110: oled_data = 16'b1111111111111111;
				14'b10110010100110: oled_data = 16'b1111111111111111;
				14'b10110100100110: oled_data = 16'b1111111111111111;
				14'b10110110100110: oled_data = 16'b1111111111111111;
				14'b10111000100110: oled_data = 16'b1111111111111111;
				14'b10111010100110: oled_data = 16'b1111111111111111;
				14'b10111100100110: oled_data = 16'b1111111111111111;
				14'b10111110100110: oled_data = 16'b1111111111111111;
				14'b00000000100111: oled_data = 16'b1111111111111111;
				14'b00000010100111: oled_data = 16'b1111111111111111;
				14'b00000100100111: oled_data = 16'b1111111111111111;
				14'b00000110100111: oled_data = 16'b1111111111111111;
				14'b00001000100111: oled_data = 16'b1111111111111111;
				14'b00001010100111: oled_data = 16'b1111111111111111;
				14'b00001100100111: oled_data = 16'b1111111111111111;
				14'b00001110100111: oled_data = 16'b1111111111111111;
				14'b00010000100111: oled_data = 16'b1111111111111111;
				14'b00010010100111: oled_data = 16'b1111111111111111;
				14'b00010100100111: oled_data = 16'b1111111111111111;
				14'b00010110100111: oled_data = 16'b1111111111111111;
				14'b00011000100111: oled_data = 16'b1111111111111111;
				14'b00011010100111: oled_data = 16'b1111111111111111;
				14'b00011100100111: oled_data = 16'b1111111111111111;
				14'b00011110100111: oled_data = 16'b1111111111111111;
				14'b00100000100111: oled_data = 16'b1111111111111111;
				14'b00100010100111: oled_data = 16'b1111111111111111;
				14'b00100100100111: oled_data = 16'b1111111111111111;
				14'b00100110100111: oled_data = 16'b1111111111111111;
				14'b00101000100111: oled_data = 16'b1111111111111111;
				14'b00101010100111: oled_data = 16'b1111111111111111;
				14'b00101100100111: oled_data = 16'b1111111111111111;
				14'b00101110100111: oled_data = 16'b1111111111111111;
				14'b00110000100111: oled_data = 16'b1111111111111111;
				14'b00110010100111: oled_data = 16'b1111111111111111;
				14'b00110100100111: oled_data = 16'b1111111111111111;
				14'b00110110100111: oled_data = 16'b1111111111111111;
				14'b00111000100111: oled_data = 16'b1111111111111111;
				14'b00111010100111: oled_data = 16'b1111111111111111;
				14'b00111100100111: oled_data = 16'b1111111111111111;
				14'b00111110100111: oled_data = 16'b1111111111111111;
				14'b01000000100111: oled_data = 16'b1111111111111111;
				14'b01000010100111: oled_data = 16'b1111111111111111;
				14'b01000100100111: oled_data = 16'b1111111111111111;
				14'b01000110100111: oled_data = 16'b1111111111111111;
				14'b01001000100111: oled_data = 16'b1111111111111111;
				14'b01001010100111: oled_data = 16'b1111111111111111;
				14'b01001100100111: oled_data = 16'b1111111111111111;
				14'b01001110100111: oled_data = 16'b1111111111111111;
				14'b01010000100111: oled_data = 16'b1111111111111111;
				14'b01010010100111: oled_data = 16'b1111111111111111;
				14'b01010100100111: oled_data = 16'b1111111111111111;
				14'b01010110100111: oled_data = 16'b1111111111111111;
				14'b01011000100111: oled_data = 16'b1111111111111111;
				14'b01011010100111: oled_data = 16'b1111111111111111;
				14'b01011100100111: oled_data = 16'b1111111111111111;
				14'b01011110100111: oled_data = 16'b1111111111111111;
				14'b01100000100111: oled_data = 16'b1111111111111111;
				14'b01100010100111: oled_data = 16'b1111111111111111;
				14'b01100100100111: oled_data = 16'b1111111111111111;
				14'b01100110100111: oled_data = 16'b1111111111111111;
				14'b01101000100111: oled_data = 16'b1111111111111111;
				14'b01101010100111: oled_data = 16'b1111111111111111;
				14'b01101100100111: oled_data = 16'b1111111111111111;
				14'b01101110100111: oled_data = 16'b1111111111111111;
				14'b01110000100111: oled_data = 16'b1111111111111111;
				14'b01110010100111: oled_data = 16'b1111111111111111;
				14'b01110100100111: oled_data = 16'b1111111111111111;
				14'b01110110100111: oled_data = 16'b1111111111111111;
				14'b01111000100111: oled_data = 16'b1111111111111111;
				14'b01111010100111: oled_data = 16'b1111111111111111;
				14'b01111100100111: oled_data = 16'b1111111111111111;
				14'b01111110100111: oled_data = 16'b1111111111111111;
				14'b10000000100111: oled_data = 16'b1111111111111111;
				14'b10000010100111: oled_data = 16'b1111111111111111;
				14'b10000100100111: oled_data = 16'b1111111111111111;
				14'b10000110100111: oled_data = 16'b1111111111111111;
				14'b10001000100111: oled_data = 16'b1111111111111111;
				14'b10001010100111: oled_data = 16'b1111111111111111;
				14'b10001100100111: oled_data = 16'b1111111111111111;
				14'b10001110100111: oled_data = 16'b1111111111111111;
				14'b10010000100111: oled_data = 16'b1111111111111111;
				14'b10010010100111: oled_data = 16'b1111111111111111;
				14'b10010100100111: oled_data = 16'b1111111111111111;
				14'b10010110100111: oled_data = 16'b1111111111111111;
				14'b10011000100111: oled_data = 16'b1111111111111111;
				14'b10011010100111: oled_data = 16'b1111111111111111;
				14'b10011100100111: oled_data = 16'b1111111111111111;
				14'b10011110100111: oled_data = 16'b1111111111111111;
				14'b10100000100111: oled_data = 16'b1111111111111111;
				14'b10100010100111: oled_data = 16'b1111111111111111;
				14'b10100100100111: oled_data = 16'b1111111111111111;
				14'b10100110100111: oled_data = 16'b1111111111111111;
				14'b10101000100111: oled_data = 16'b1111111111111111;
				14'b10101010100111: oled_data = 16'b1111111111111111;
				14'b10101100100111: oled_data = 16'b1111111111111111;
				14'b10101110100111: oled_data = 16'b1111111111111111;
				14'b10110000100111: oled_data = 16'b1111111111111111;
				14'b10110010100111: oled_data = 16'b1111111111111111;
				14'b10110100100111: oled_data = 16'b1111111111111111;
				14'b10110110100111: oled_data = 16'b1111111111111111;
				14'b10111000100111: oled_data = 16'b1111111111111111;
				14'b10111010100111: oled_data = 16'b1111111111111111;
				14'b10111100100111: oled_data = 16'b1111111111111111;
				14'b10111110100111: oled_data = 16'b1111111111111111;
				14'b00000000101000: oled_data = 16'b1111111111111111;
				14'b00000010101000: oled_data = 16'b1111111111111111;
				14'b00000100101000: oled_data = 16'b1111111111111111;
				14'b00000110101000: oled_data = 16'b1111111111111111;
				14'b00001000101000: oled_data = 16'b1111111111111111;
				14'b00001010101000: oled_data = 16'b1111111111111111;
				14'b00001100101000: oled_data = 16'b1111111111111111;
				14'b00001110101000: oled_data = 16'b1111111111111111;
				14'b00010000101000: oled_data = 16'b1111111111111111;
				14'b00010010101000: oled_data = 16'b1111111111111111;
				14'b00010100101000: oled_data = 16'b1111111111111111;
				14'b00010110101000: oled_data = 16'b1111111111111111;
				14'b00011000101000: oled_data = 16'b1111111111111111;
				14'b00011010101000: oled_data = 16'b1111111111111111;
				14'b00011100101000: oled_data = 16'b1111111111111111;
				14'b00011110101000: oled_data = 16'b1111111111111111;
				14'b00100000101000: oled_data = 16'b1111111111111111;
				14'b00100010101000: oled_data = 16'b1111111111111111;
				14'b00100100101000: oled_data = 16'b1111111111111111;
				14'b00100110101000: oled_data = 16'b1111111111111111;
				14'b00101000101000: oled_data = 16'b1111111111111111;
				14'b00101010101000: oled_data = 16'b1111111111111111;
				14'b00101100101000: oled_data = 16'b1111111111111111;
				14'b00101110101000: oled_data = 16'b1111111111111111;
				14'b00110000101000: oled_data = 16'b1111111111111111;
				14'b00110010101000: oled_data = 16'b1111111111111111;
				14'b00110100101000: oled_data = 16'b1111111111111111;
				14'b00110110101000: oled_data = 16'b1111111111111111;
				14'b00111000101000: oled_data = 16'b1111111111111111;
				14'b00111010101000: oled_data = 16'b1111111111111111;
				14'b00111100101000: oled_data = 16'b1111111111111111;
				14'b00111110101000: oled_data = 16'b1111111111111111;
				14'b01000000101000: oled_data = 16'b1111111111111111;
				14'b01000010101000: oled_data = 16'b1111111111111111;
				14'b01000100101000: oled_data = 16'b1111111111111111;
				14'b01000110101000: oled_data = 16'b1111111111111111;
				14'b01001000101000: oled_data = 16'b1111111111111111;
				14'b01001010101000: oled_data = 16'b1111111111111111;
				14'b01001100101000: oled_data = 16'b1111111111111111;
				14'b01001110101000: oled_data = 16'b1111111111111111;
				14'b01010000101000: oled_data = 16'b1111111111111111;
				14'b01010010101000: oled_data = 16'b1111111111111111;
				14'b01010100101000: oled_data = 16'b1111111111111111;
				14'b01010110101000: oled_data = 16'b1111111111111111;
				14'b01011000101000: oled_data = 16'b1111111111111111;
				14'b01011010101000: oled_data = 16'b1111111111111111;
				14'b01011100101000: oled_data = 16'b1111111111111111;
				14'b01011110101000: oled_data = 16'b1111111111111111;
				14'b01100000101000: oled_data = 16'b1111111111111111;
				14'b01100010101000: oled_data = 16'b1111111111111111;
				14'b01100100101000: oled_data = 16'b1111111111111111;
				14'b01100110101000: oled_data = 16'b1111111111111111;
				14'b01101000101000: oled_data = 16'b1111111111111111;
				14'b01101010101000: oled_data = 16'b1111111111111111;
				14'b01101100101000: oled_data = 16'b1111111111111111;
				14'b01101110101000: oled_data = 16'b1111111111111111;
				14'b01110000101000: oled_data = 16'b1111111111111111;
				14'b01110010101000: oled_data = 16'b1111111111111111;
				14'b01110100101000: oled_data = 16'b1111111111111111;
				14'b01110110101000: oled_data = 16'b1111111111111111;
				14'b01111000101000: oled_data = 16'b1111111111111111;
				14'b01111010101000: oled_data = 16'b1111111111111111;
				14'b01111100101000: oled_data = 16'b1111111111111111;
				14'b01111110101000: oled_data = 16'b1111111111111111;
				14'b10000000101000: oled_data = 16'b1111111111111111;
				14'b10000010101000: oled_data = 16'b1111111111111111;
				14'b10000100101000: oled_data = 16'b1111111111111111;
				14'b10000110101000: oled_data = 16'b1111111111111111;
				14'b10001000101000: oled_data = 16'b1111111111111111;
				14'b10001010101000: oled_data = 16'b1111111111111111;
				14'b10001100101000: oled_data = 16'b1111111111111111;
				14'b10001110101000: oled_data = 16'b1111111111111111;
				14'b10010000101000: oled_data = 16'b1111111111111111;
				14'b10010010101000: oled_data = 16'b1111111111111111;
				14'b10010100101000: oled_data = 16'b1111111111111111;
				14'b10010110101000: oled_data = 16'b1111111111111111;
				14'b10011000101000: oled_data = 16'b1111111111111111;
				14'b10011010101000: oled_data = 16'b1111111111111111;
				14'b10011100101000: oled_data = 16'b1111111111111111;
				14'b10011110101000: oled_data = 16'b1111111111111111;
				14'b10100000101000: oled_data = 16'b1111111111111111;
				14'b10100010101000: oled_data = 16'b1111111111111111;
				14'b10100100101000: oled_data = 16'b1111111111111111;
				14'b10100110101000: oled_data = 16'b1111111111111111;
				14'b10101000101000: oled_data = 16'b1111111111111111;
				14'b10101010101000: oled_data = 16'b1111111111111111;
				14'b10101100101000: oled_data = 16'b1111111111111111;
				14'b10101110101000: oled_data = 16'b1111111111111111;
				14'b10110000101000: oled_data = 16'b1111111111111111;
				14'b10110010101000: oled_data = 16'b1111111111111111;
				14'b10110100101000: oled_data = 16'b1111111111111111;
				14'b10110110101000: oled_data = 16'b1111111111111111;
				14'b10111000101000: oled_data = 16'b1111111111111111;
				14'b10111010101000: oled_data = 16'b1111111111111111;
				14'b10111100101000: oled_data = 16'b1111111111111111;
				14'b10111110101000: oled_data = 16'b1111111111111111;
				14'b00000000101001: oled_data = 16'b1111111111111111;
				14'b00000010101001: oled_data = 16'b1111111111111111;
				14'b00000100101001: oled_data = 16'b1111111111111111;
				14'b00000110101001: oled_data = 16'b1111111111111111;
				14'b00001000101001: oled_data = 16'b1111111111111111;
				14'b00001010101001: oled_data = 16'b1111111111111111;
				14'b00001100101001: oled_data = 16'b1111111111111111;
				14'b00001110101001: oled_data = 16'b1111111111111111;
				14'b00010000101001: oled_data = 16'b1111111111111111;
				14'b00010010101001: oled_data = 16'b1111111111111111;
				14'b00010100101001: oled_data = 16'b1111111111111111;
				14'b00010110101001: oled_data = 16'b1111111111111111;
				14'b00011000101001: oled_data = 16'b1111111111111111;
				14'b00011010101001: oled_data = 16'b1111111111111111;
				14'b00011100101001: oled_data = 16'b1111111111111111;
				14'b00011110101001: oled_data = 16'b1111111111111111;
				14'b00100000101001: oled_data = 16'b1111111111111111;
				14'b00100010101001: oled_data = 16'b1111111111111111;
				14'b00100100101001: oled_data = 16'b1111111111111111;
				14'b00100110101001: oled_data = 16'b1111111111111111;
				14'b00101000101001: oled_data = 16'b1111111111111111;
				14'b00101010101001: oled_data = 16'b1111111111111111;
				14'b00101100101001: oled_data = 16'b1111111111111111;
				14'b00101110101001: oled_data = 16'b1111111111111111;
				14'b00110000101001: oled_data = 16'b1111111111111111;
				14'b00110010101001: oled_data = 16'b1111111111111111;
				14'b00110100101001: oled_data = 16'b1111111111111111;
				14'b00110110101001: oled_data = 16'b1111111111111111;
				14'b00111000101001: oled_data = 16'b1111111111111111;
				14'b00111010101001: oled_data = 16'b1111111111111111;
				14'b00111100101001: oled_data = 16'b1111111111111111;
				14'b00111110101001: oled_data = 16'b1111111111111111;
				14'b01000000101001: oled_data = 16'b1111111111111111;
				14'b01000010101001: oled_data = 16'b1111111111111111;
				14'b01000100101001: oled_data = 16'b1111111111111111;
				14'b01000110101001: oled_data = 16'b1111111111111111;
				14'b01001000101001: oled_data = 16'b1111111111111111;
				14'b01001010101001: oled_data = 16'b1111111111111111;
				14'b01001100101001: oled_data = 16'b1111111111111111;
				14'b01001110101001: oled_data = 16'b1111111111111111;
				14'b01010000101001: oled_data = 16'b1111111111111111;
				14'b01010010101001: oled_data = 16'b1111111111111111;
				14'b01010100101001: oled_data = 16'b1111111111111111;
				14'b01010110101001: oled_data = 16'b1111111111111111;
				14'b01011000101001: oled_data = 16'b1111111111111111;
				14'b01011010101001: oled_data = 16'b1111111111111111;
				14'b01011100101001: oled_data = 16'b1111111111111111;
				14'b01011110101001: oled_data = 16'b1111111111111111;
				14'b01100000101001: oled_data = 16'b1111111111111111;
				14'b01100010101001: oled_data = 16'b1111111111111111;
				14'b01100100101001: oled_data = 16'b1111111111111111;
				14'b01100110101001: oled_data = 16'b1111111111111111;
				14'b01101000101001: oled_data = 16'b1111111111111111;
				14'b01101010101001: oled_data = 16'b1111111111111111;
				14'b01101100101001: oled_data = 16'b1111111111111111;
				14'b01101110101001: oled_data = 16'b1111111111111111;
				14'b01110000101001: oled_data = 16'b1111111111111111;
				14'b01110010101001: oled_data = 16'b1111111111111111;
				14'b01110100101001: oled_data = 16'b1111111111111111;
				14'b01110110101001: oled_data = 16'b1111111111111111;
				14'b01111000101001: oled_data = 16'b1111111111111111;
				14'b01111010101001: oled_data = 16'b1111111111111111;
				14'b01111100101001: oled_data = 16'b1111111111111111;
				14'b01111110101001: oled_data = 16'b1111111111111111;
				14'b10000000101001: oled_data = 16'b1111111111111111;
				14'b10000010101001: oled_data = 16'b1111111111111111;
				14'b10000100101001: oled_data = 16'b1111111111111111;
				14'b10000110101001: oled_data = 16'b1111111111111111;
				14'b10001000101001: oled_data = 16'b1111111111111111;
				14'b10001010101001: oled_data = 16'b1111111111111111;
				14'b10001100101001: oled_data = 16'b1111111111111111;
				14'b10001110101001: oled_data = 16'b1111111111111111;
				14'b10010000101001: oled_data = 16'b1111111111111111;
				14'b10010010101001: oled_data = 16'b1111111111111111;
				14'b10010100101001: oled_data = 16'b1111111111111111;
				14'b10010110101001: oled_data = 16'b1111111111111111;
				14'b10011000101001: oled_data = 16'b1111111111111111;
				14'b10011010101001: oled_data = 16'b1111111111111111;
				14'b10011100101001: oled_data = 16'b1111111111111111;
				14'b10011110101001: oled_data = 16'b1111111111111111;
				14'b10100000101001: oled_data = 16'b1111111111111111;
				14'b10100010101001: oled_data = 16'b1111111111111111;
				14'b10100100101001: oled_data = 16'b1111111111111111;
				14'b10100110101001: oled_data = 16'b1111111111111111;
				14'b10101000101001: oled_data = 16'b1111111111111111;
				14'b10101010101001: oled_data = 16'b1111111111111111;
				14'b10101100101001: oled_data = 16'b1111111111111111;
				14'b10101110101001: oled_data = 16'b1111111111111111;
				14'b10110000101001: oled_data = 16'b1111111111111111;
				14'b10110010101001: oled_data = 16'b1111111111111111;
				14'b10110100101001: oled_data = 16'b1111111111111111;
				14'b10110110101001: oled_data = 16'b1111111111111111;
				14'b10111000101001: oled_data = 16'b1111111111111111;
				14'b10111010101001: oled_data = 16'b1111111111111111;
				14'b10111100101001: oled_data = 16'b1111111111111111;
				14'b10111110101001: oled_data = 16'b1111111111111111;
				14'b00000000101010: oled_data = 16'b1111111111111111;
				14'b00000010101010: oled_data = 16'b1111111111111111;
				14'b00000100101010: oled_data = 16'b1111111111111111;
				14'b00000110101010: oled_data = 16'b1111111111111111;
				14'b00001000101010: oled_data = 16'b1111111111111111;
				14'b00001010101010: oled_data = 16'b1111111111111111;
				14'b00001100101010: oled_data = 16'b1111111111111111;
				14'b00001110101010: oled_data = 16'b1111111111111111;
				14'b00010000101010: oled_data = 16'b1111111111111111;
				14'b00010010101010: oled_data = 16'b1111111111111111;
				14'b00010100101010: oled_data = 16'b1111111111111111;
				14'b00010110101010: oled_data = 16'b1111111111111111;
				14'b00011000101010: oled_data = 16'b1111111111111111;
				14'b00011010101010: oled_data = 16'b1111111111111111;
				14'b00011100101010: oled_data = 16'b1111111111111111;
				14'b00011110101010: oled_data = 16'b1111111111111111;
				14'b00100000101010: oled_data = 16'b1111111111111111;
				14'b00100010101010: oled_data = 16'b1111111111111111;
				14'b00100100101010: oled_data = 16'b1111111111111111;
				14'b00100110101010: oled_data = 16'b1111111111111111;
				14'b00101000101010: oled_data = 16'b1111111111111111;
				14'b00101010101010: oled_data = 16'b1111111111111111;
				14'b00101100101010: oled_data = 16'b1111111111111111;
				14'b00101110101010: oled_data = 16'b1111111111111111;
				14'b00110000101010: oled_data = 16'b1111111111111111;
				14'b00110010101010: oled_data = 16'b1111111111111111;
				14'b00110100101010: oled_data = 16'b1111111111111111;
				14'b00110110101010: oled_data = 16'b1111111111111111;
				14'b00111000101010: oled_data = 16'b1111111111111111;
				14'b00111010101010: oled_data = 16'b1111111111111111;
				14'b00111100101010: oled_data = 16'b1111111111111111;
				14'b00111110101010: oled_data = 16'b1111111111111111;
				14'b01000000101010: oled_data = 16'b1111111111111111;
				14'b01000010101010: oled_data = 16'b1111111111111111;
				14'b01000100101010: oled_data = 16'b1111111111111111;
				14'b01000110101010: oled_data = 16'b1111111111111111;
				14'b01001000101010: oled_data = 16'b1111111111111111;
				14'b01001010101010: oled_data = 16'b1111111111111111;
				14'b01001100101010: oled_data = 16'b1111111111111111;
				14'b01001110101010: oled_data = 16'b1111111111111111;
				14'b01010000101010: oled_data = 16'b1111111111111111;
				14'b01010010101010: oled_data = 16'b1111111111111111;
				14'b01010100101010: oled_data = 16'b1111111111111111;
				14'b01010110101010: oled_data = 16'b1111111111111111;
				14'b01011000101010: oled_data = 16'b1111111111111111;
				14'b01011010101010: oled_data = 16'b1111111111111111;
				14'b01011100101010: oled_data = 16'b1111111111111111;
				14'b01011110101010: oled_data = 16'b1111111111111111;
				14'b01100000101010: oled_data = 16'b1111111111111111;
				14'b01100010101010: oled_data = 16'b1111111111111111;
				14'b01100100101010: oled_data = 16'b1111111111111111;
				14'b01100110101010: oled_data = 16'b1111111111111111;
				14'b01101000101010: oled_data = 16'b1111111111111111;
				14'b01101010101010: oled_data = 16'b1111111111111111;
				14'b01101100101010: oled_data = 16'b1111111111111111;
				14'b01101110101010: oled_data = 16'b1111111111111111;
				14'b01110000101010: oled_data = 16'b1111111111111111;
				14'b01110010101010: oled_data = 16'b1111111111111111;
				14'b01110100101010: oled_data = 16'b1111111111111111;
				14'b01110110101010: oled_data = 16'b1111111111111111;
				14'b01111000101010: oled_data = 16'b1111111111111111;
				14'b01111010101010: oled_data = 16'b1111111111111111;
				14'b01111100101010: oled_data = 16'b1111111111111111;
				14'b01111110101010: oled_data = 16'b1111111111111111;
				14'b10000000101010: oled_data = 16'b1111111111111111;
				14'b10000010101010: oled_data = 16'b1111111111111111;
				14'b10000100101010: oled_data = 16'b1111111111111111;
				14'b10000110101010: oled_data = 16'b1111111111111111;
				14'b10001000101010: oled_data = 16'b1111111111111111;
				14'b10001010101010: oled_data = 16'b1111111111111111;
				14'b10001100101010: oled_data = 16'b1111111111111111;
				14'b10001110101010: oled_data = 16'b1111111111111111;
				14'b10010000101010: oled_data = 16'b1111111111111111;
				14'b10010010101010: oled_data = 16'b1111111111111111;
				14'b10010100101010: oled_data = 16'b1111111111111111;
				14'b10010110101010: oled_data = 16'b1111111111111111;
				14'b10011000101010: oled_data = 16'b1111111111111111;
				14'b10011010101010: oled_data = 16'b1111111111111111;
				14'b10011100101010: oled_data = 16'b1111111111111111;
				14'b10011110101010: oled_data = 16'b1111111111111111;
				14'b10100000101010: oled_data = 16'b1111111111111111;
				14'b10100010101010: oled_data = 16'b1111111111111111;
				14'b10100100101010: oled_data = 16'b1111111111111111;
				14'b10100110101010: oled_data = 16'b1111111111111111;
				14'b10101000101010: oled_data = 16'b1111111111111111;
				14'b10101010101010: oled_data = 16'b1111111111111111;
				14'b10101100101010: oled_data = 16'b1111111111111111;
				14'b10101110101010: oled_data = 16'b1111111111111111;
				14'b10110000101010: oled_data = 16'b1111111111111111;
				14'b10110010101010: oled_data = 16'b1111111111111111;
				14'b10110100101010: oled_data = 16'b1111111111111111;
				14'b10110110101010: oled_data = 16'b1111111111111111;
				14'b10111000101010: oled_data = 16'b1111111111111111;
				14'b10111010101010: oled_data = 16'b1111111111111111;
				14'b10111100101010: oled_data = 16'b1111111111111111;
				14'b10111110101010: oled_data = 16'b1111111111111111;
				14'b00000000101011: oled_data = 16'b1111111111111111;
				14'b00000010101011: oled_data = 16'b1111111111111111;
				14'b00000100101011: oled_data = 16'b1111111111111111;
				14'b00000110101011: oled_data = 16'b1111111111111111;
				14'b00001000101011: oled_data = 16'b1111111111111111;
				14'b00001010101011: oled_data = 16'b1111111111111111;
				14'b00001100101011: oled_data = 16'b1111111111111111;
				14'b00001110101011: oled_data = 16'b1111111111111111;
				14'b00010000101011: oled_data = 16'b1111111111111111;
				14'b00010010101011: oled_data = 16'b1111111111111111;
				14'b00010100101011: oled_data = 16'b1111111111111111;
				14'b00010110101011: oled_data = 16'b1111111111111111;
				14'b00011000101011: oled_data = 16'b1111111111111111;
				14'b00011010101011: oled_data = 16'b1111111111111111;
				14'b00011100101011: oled_data = 16'b1111111111111111;
				14'b00011110101011: oled_data = 16'b1111111111111111;
				14'b00100000101011: oled_data = 16'b1111111111111111;
				14'b00100010101011: oled_data = 16'b1111111111111111;
				14'b00100100101011: oled_data = 16'b1111111111111111;
				14'b00100110101011: oled_data = 16'b1111111111111111;
				14'b00101000101011: oled_data = 16'b1111111111111111;
				14'b00101010101011: oled_data = 16'b1111111111111111;
				14'b00101100101011: oled_data = 16'b1111111111111111;
				14'b00101110101011: oled_data = 16'b1111111111111111;
				14'b00110000101011: oled_data = 16'b1111111111111111;
				14'b00110010101011: oled_data = 16'b1111111111111111;
				14'b00110100101011: oled_data = 16'b1111111111111111;
				14'b00110110101011: oled_data = 16'b1111111111111111;
				14'b00111000101011: oled_data = 16'b1111111111111111;
				14'b00111010101011: oled_data = 16'b1111111111111111;
				14'b00111100101011: oled_data = 16'b1111111111111111;
				14'b00111110101011: oled_data = 16'b1111111111111111;
				14'b01000000101011: oled_data = 16'b1111111111111111;
				14'b01000010101011: oled_data = 16'b1111111111111111;
				14'b01000100101011: oled_data = 16'b1111111111111111;
				14'b01000110101011: oled_data = 16'b1111111111111111;
				14'b01001000101011: oled_data = 16'b1111111111111111;
				14'b01001010101011: oled_data = 16'b1111111111111111;
				14'b01001100101011: oled_data = 16'b1111111111111111;
				14'b01001110101011: oled_data = 16'b1111111111111111;
				14'b01010000101011: oled_data = 16'b1111111111111111;
				14'b01010010101011: oled_data = 16'b1111111111111111;
				14'b01010100101011: oled_data = 16'b1111111111111111;
				14'b01010110101011: oled_data = 16'b1111111111111111;
				14'b01011000101011: oled_data = 16'b1111111111111111;
				14'b01011010101011: oled_data = 16'b1111111111111111;
				14'b01011100101011: oled_data = 16'b1111111111111111;
				14'b01011110101011: oled_data = 16'b1111111111111111;
				14'b01100000101011: oled_data = 16'b1111111111111111;
				14'b01100010101011: oled_data = 16'b1111111111111111;
				14'b01100100101011: oled_data = 16'b1111111111111111;
				14'b01100110101011: oled_data = 16'b1111111111111111;
				14'b01101000101011: oled_data = 16'b1111111111111111;
				14'b01101010101011: oled_data = 16'b1111111111111111;
				14'b01101100101011: oled_data = 16'b1111111111111111;
				14'b01101110101011: oled_data = 16'b1111111111111111;
				14'b01110000101011: oled_data = 16'b1111111111111111;
				14'b01110010101011: oled_data = 16'b1111111111111111;
				14'b01110100101011: oled_data = 16'b1111111111111111;
				14'b01110110101011: oled_data = 16'b1111111111111111;
				14'b01111000101011: oled_data = 16'b1111111111111111;
				14'b01111010101011: oled_data = 16'b1111111111111111;
				14'b01111100101011: oled_data = 16'b1111111111111111;
				14'b01111110101011: oled_data = 16'b1111111111111111;
				14'b10000000101011: oled_data = 16'b1111111111111111;
				14'b10000010101011: oled_data = 16'b1111111111111111;
				14'b10000100101011: oled_data = 16'b1111111111111111;
				14'b10000110101011: oled_data = 16'b1111111111111111;
				14'b10001000101011: oled_data = 16'b1111111111111111;
				14'b10001010101011: oled_data = 16'b1111111111111111;
				14'b10001100101011: oled_data = 16'b1111111111111111;
				14'b10001110101011: oled_data = 16'b1111111111111111;
				14'b10010000101011: oled_data = 16'b1111111111111111;
				14'b10010010101011: oled_data = 16'b1111111111111111;
				14'b10010100101011: oled_data = 16'b1111111111111111;
				14'b10010110101011: oled_data = 16'b1111111111111111;
				14'b10011000101011: oled_data = 16'b1111111111111111;
				14'b10011010101011: oled_data = 16'b1111111111111111;
				14'b10011100101011: oled_data = 16'b1111111111111111;
				14'b10011110101011: oled_data = 16'b1111111111111111;
				14'b10100000101011: oled_data = 16'b1111111111111111;
				14'b10100010101011: oled_data = 16'b1111111111111111;
				14'b10100100101011: oled_data = 16'b1111111111111111;
				14'b10100110101011: oled_data = 16'b1111111111111111;
				14'b10101000101011: oled_data = 16'b1111111111111111;
				14'b10101010101011: oled_data = 16'b1111111111111111;
				14'b10101100101011: oled_data = 16'b1111111111111111;
				14'b10101110101011: oled_data = 16'b1111111111111111;
				14'b10110000101011: oled_data = 16'b1111111111111111;
				14'b10110010101011: oled_data = 16'b1111111111111111;
				14'b10110100101011: oled_data = 16'b1111111111111111;
				14'b10110110101011: oled_data = 16'b1111111111111111;
				14'b10111000101011: oled_data = 16'b1111111111111111;
				14'b10111010101011: oled_data = 16'b1111111111111111;
				14'b10111100101011: oled_data = 16'b1111111111111111;
				14'b10111110101011: oled_data = 16'b1111111111111111;
				14'b00000000101100: oled_data = 16'b1111111111111111;
				14'b00000010101100: oled_data = 16'b1111111111111111;
				14'b00000100101100: oled_data = 16'b1111111111111111;
				14'b00000110101100: oled_data = 16'b1111111111111111;
				14'b00001000101100: oled_data = 16'b1111111111111111;
				14'b00001010101100: oled_data = 16'b1111111111111111;
				14'b00001100101100: oled_data = 16'b1111111111111111;
				14'b00001110101100: oled_data = 16'b1111111111111111;
				14'b00010000101100: oled_data = 16'b1111111111111111;
				14'b00010010101100: oled_data = 16'b1111111111111111;
				14'b00010100101100: oled_data = 16'b1111111111111111;
				14'b00010110101100: oled_data = 16'b1111111111111111;
				14'b00011000101100: oled_data = 16'b1111111111111111;
				14'b00011010101100: oled_data = 16'b1111111111111111;
				14'b00011100101100: oled_data = 16'b1111111111111111;
				14'b00011110101100: oled_data = 16'b1111111111111111;
				14'b00100000101100: oled_data = 16'b1111111111111111;
				14'b00100010101100: oled_data = 16'b1111111111111111;
				14'b00100100101100: oled_data = 16'b1111111111111111;
				14'b00100110101100: oled_data = 16'b1111111111111111;
				14'b00101000101100: oled_data = 16'b1111111111111111;
				14'b00101010101100: oled_data = 16'b1111111111111111;
				14'b00101100101100: oled_data = 16'b1111111111111111;
				14'b00101110101100: oled_data = 16'b1111111111111111;
				14'b00110000101100: oled_data = 16'b1111111111111111;
				14'b00110010101100: oled_data = 16'b1111111111111111;
				14'b00110100101100: oled_data = 16'b1111111111111111;
				14'b00110110101100: oled_data = 16'b1111111111111111;
				14'b00111000101100: oled_data = 16'b1111111111111111;
				14'b00111010101100: oled_data = 16'b1111111111111111;
				14'b00111100101100: oled_data = 16'b1111111111111111;
				14'b00111110101100: oled_data = 16'b1111111111111111;
				14'b01000000101100: oled_data = 16'b1111111111111111;
				14'b01000010101100: oled_data = 16'b1111111111111111;
				14'b01000100101100: oled_data = 16'b1111111111111111;
				14'b01000110101100: oled_data = 16'b1111111111111111;
				14'b01001000101100: oled_data = 16'b1111111111111111;
				14'b01001010101100: oled_data = 16'b1111111111111111;
				14'b01001100101100: oled_data = 16'b1111111111111111;
				14'b01001110101100: oled_data = 16'b1111111111111111;
				14'b01010000101100: oled_data = 16'b1111111111111111;
				14'b01010010101100: oled_data = 16'b1111111111111111;
				14'b01010100101100: oled_data = 16'b1111111111111111;
				14'b01010110101100: oled_data = 16'b1111111111111111;
				14'b01011000101100: oled_data = 16'b1111111111111111;
				14'b01011010101100: oled_data = 16'b1111111111111111;
				14'b01011100101100: oled_data = 16'b1111111111111111;
				14'b01011110101100: oled_data = 16'b1111111111111111;
				14'b01100000101100: oled_data = 16'b1111111111111111;
				14'b01100010101100: oled_data = 16'b1111111111111111;
				14'b01100100101100: oled_data = 16'b1111111111111111;
				14'b01100110101100: oled_data = 16'b1111111111111111;
				14'b01101000101100: oled_data = 16'b1111111111111111;
				14'b01101010101100: oled_data = 16'b1111111111111111;
				14'b01101100101100: oled_data = 16'b1111111111111111;
				14'b01101110101100: oled_data = 16'b1111111111111111;
				14'b01110000101100: oled_data = 16'b1111111111111111;
				14'b01110010101100: oled_data = 16'b1111111111111111;
				14'b01110100101100: oled_data = 16'b1111111111111111;
				14'b01110110101100: oled_data = 16'b1111111111111111;
				14'b01111000101100: oled_data = 16'b1111111111111111;
				14'b01111010101100: oled_data = 16'b1111111111111111;
				14'b01111100101100: oled_data = 16'b1111111111111111;
				14'b01111110101100: oled_data = 16'b1111111111111111;
				14'b10000000101100: oled_data = 16'b1111111111111111;
				14'b10000010101100: oled_data = 16'b1111111111111111;
				14'b10000100101100: oled_data = 16'b1111111111111111;
				14'b10000110101100: oled_data = 16'b1111111111111111;
				14'b10001000101100: oled_data = 16'b1111111111111111;
				14'b10001010101100: oled_data = 16'b1111111111111111;
				14'b10001100101100: oled_data = 16'b1111111111111111;
				14'b10001110101100: oled_data = 16'b1111111111111111;
				14'b10010000101100: oled_data = 16'b1111111111111111;
				14'b10010010101100: oled_data = 16'b1111111111111111;
				14'b10010100101100: oled_data = 16'b1111111111111111;
				14'b10010110101100: oled_data = 16'b1111111111111111;
				14'b10011000101100: oled_data = 16'b1111111111111111;
				14'b10011010101100: oled_data = 16'b1111111111111111;
				14'b10011100101100: oled_data = 16'b1111111111111111;
				14'b10011110101100: oled_data = 16'b1111111111111111;
				14'b10100000101100: oled_data = 16'b1111111111111111;
				14'b10100010101100: oled_data = 16'b1111111111111111;
				14'b10100100101100: oled_data = 16'b1111111111111111;
				14'b10100110101100: oled_data = 16'b1111111111111111;
				14'b10101000101100: oled_data = 16'b1111111111111111;
				14'b10101010101100: oled_data = 16'b1111111111111111;
				14'b10101100101100: oled_data = 16'b1111111111111111;
				14'b10101110101100: oled_data = 16'b1111111111111111;
				14'b10110000101100: oled_data = 16'b1111111111111111;
				14'b10110010101100: oled_data = 16'b1111111111111111;
				14'b10110100101100: oled_data = 16'b1111111111111111;
				14'b10110110101100: oled_data = 16'b1111111111111111;
				14'b10111000101100: oled_data = 16'b1111111111111111;
				14'b10111010101100: oled_data = 16'b1111111111111111;
				14'b10111100101100: oled_data = 16'b1111111111111111;
				14'b10111110101100: oled_data = 16'b1111111111111111;
				14'b00000000101101: oled_data = 16'b1111111111111111;
				14'b00000010101101: oled_data = 16'b1111111111111111;
				14'b00000100101101: oled_data = 16'b1111111111111111;
				14'b00000110101101: oled_data = 16'b1111111111111111;
				14'b00001000101101: oled_data = 16'b1111111111111111;
				14'b00001010101101: oled_data = 16'b1111111111111111;
				14'b00001100101101: oled_data = 16'b1111111111111111;
				14'b00001110101101: oled_data = 16'b1111111111111111;
				14'b00010000101101: oled_data = 16'b1111111111111111;
				14'b00010010101101: oled_data = 16'b1111111111111111;
				14'b00010100101101: oled_data = 16'b1111111111111111;
				14'b00010110101101: oled_data = 16'b1111111111111111;
				14'b00011000101101: oled_data = 16'b1111111111111111;
				14'b00011010101101: oled_data = 16'b1111111111111111;
				14'b00011100101101: oled_data = 16'b1111111111111111;
				14'b00011110101101: oled_data = 16'b1111111111111111;
				14'b00100000101101: oled_data = 16'b1111111111111111;
				14'b00100010101101: oled_data = 16'b1111111111111111;
				14'b00100100101101: oled_data = 16'b1111111111111111;
				14'b00100110101101: oled_data = 16'b1111111111111111;
				14'b00101000101101: oled_data = 16'b1111111111111111;
				14'b00101010101101: oled_data = 16'b1111111111111111;
				14'b00101100101101: oled_data = 16'b1111111111111111;
				14'b00101110101101: oled_data = 16'b1111111111111111;
				14'b00110000101101: oled_data = 16'b1111111111111111;
				14'b00110010101101: oled_data = 16'b1111111111111111;
				14'b00110100101101: oled_data = 16'b1111111111111111;
				14'b00110110101101: oled_data = 16'b1111111111111111;
				14'b00111000101101: oled_data = 16'b1111111111111111;
				14'b00111010101101: oled_data = 16'b1111111111111111;
				14'b00111100101101: oled_data = 16'b1111111111111111;
				14'b00111110101101: oled_data = 16'b1111111111111111;
				14'b01000000101101: oled_data = 16'b1111111111111111;
				14'b01000010101101: oled_data = 16'b1111111111111111;
				14'b01000100101101: oled_data = 16'b1111111111111111;
				14'b01000110101101: oled_data = 16'b1111111111111111;
				14'b01001000101101: oled_data = 16'b1111111111111111;
				14'b01001010101101: oled_data = 16'b1111111111111111;
				14'b01001100101101: oled_data = 16'b1111111111111111;
				14'b01001110101101: oled_data = 16'b1111111111111111;
				14'b01010000101101: oled_data = 16'b1111111111111111;
				14'b01010010101101: oled_data = 16'b1111111111111111;
				14'b01010100101101: oled_data = 16'b1111111111111111;
				14'b01010110101101: oled_data = 16'b1111111111111111;
				14'b01011000101101: oled_data = 16'b1111111111111111;
				14'b01011010101101: oled_data = 16'b1111111111111111;
				14'b01011100101101: oled_data = 16'b1111111111111111;
				14'b01011110101101: oled_data = 16'b1111111111111111;
				14'b01100000101101: oled_data = 16'b1111111111111111;
				14'b01100010101101: oled_data = 16'b1111111111111111;
				14'b01100100101101: oled_data = 16'b1111111111111111;
				14'b01100110101101: oled_data = 16'b1111111111111111;
				14'b01101000101101: oled_data = 16'b1111111111111111;
				14'b01101010101101: oled_data = 16'b1111111111111111;
				14'b01101100101101: oled_data = 16'b1111111111111111;
				14'b01101110101101: oled_data = 16'b1111111111111111;
				14'b01110000101101: oled_data = 16'b1111111111111111;
				14'b01110010101101: oled_data = 16'b1111111111111111;
				14'b01110100101101: oled_data = 16'b1111111111111111;
				14'b01110110101101: oled_data = 16'b1111111111111111;
				14'b01111000101101: oled_data = 16'b1111111111111111;
				14'b01111010101101: oled_data = 16'b1111111111111111;
				14'b01111100101101: oled_data = 16'b1111111111111111;
				14'b01111110101101: oled_data = 16'b1111111111111111;
				14'b10000000101101: oled_data = 16'b1111111111111111;
				14'b10000010101101: oled_data = 16'b1111111111111111;
				14'b10000100101101: oled_data = 16'b1111111111111111;
				14'b10000110101101: oled_data = 16'b1111111111111111;
				14'b10001000101101: oled_data = 16'b1111111111111111;
				14'b10001010101101: oled_data = 16'b1111111111111111;
				14'b10001100101101: oled_data = 16'b1111111111111111;
				14'b10001110101101: oled_data = 16'b1111111111111111;
				14'b10010000101101: oled_data = 16'b1111111111111111;
				14'b10010010101101: oled_data = 16'b1111111111111111;
				14'b10010100101101: oled_data = 16'b1111111111111111;
				14'b10010110101101: oled_data = 16'b1111111111111111;
				14'b10011000101101: oled_data = 16'b1111111111111111;
				14'b10011010101101: oled_data = 16'b1111111111111111;
				14'b10011100101101: oled_data = 16'b1111111111111111;
				14'b10011110101101: oled_data = 16'b1111111111111111;
				14'b10100000101101: oled_data = 16'b1111111111111111;
				14'b10100010101101: oled_data = 16'b1111111111111111;
				14'b10100100101101: oled_data = 16'b1111111111111111;
				14'b10100110101101: oled_data = 16'b1111111111111111;
				14'b10101000101101: oled_data = 16'b1111111111111111;
				14'b10101010101101: oled_data = 16'b1111111111111111;
				14'b10101100101101: oled_data = 16'b1111111111111111;
				14'b10101110101101: oled_data = 16'b1111111111111111;
				14'b10110000101101: oled_data = 16'b1111111111111111;
				14'b10110010101101: oled_data = 16'b1111111111111111;
				14'b10110100101101: oled_data = 16'b1111111111111111;
				14'b10110110101101: oled_data = 16'b1111111111111111;
				14'b10111000101101: oled_data = 16'b1111111111111111;
				14'b10111010101101: oled_data = 16'b1111111111111111;
				14'b10111100101101: oled_data = 16'b1111111111111111;
				14'b10111110101101: oled_data = 16'b1111111111111111;
				14'b00000000101110: oled_data = 16'b1111111111111111;
				14'b00000010101110: oled_data = 16'b1111111111111111;
				14'b00000100101110: oled_data = 16'b1111111111111111;
				14'b00000110101110: oled_data = 16'b1111111111111111;
				14'b00001000101110: oled_data = 16'b1111111111111111;
				14'b00001010101110: oled_data = 16'b1111111111111111;
				14'b00001100101110: oled_data = 16'b1111111111111111;
				14'b00001110101110: oled_data = 16'b1111111111111111;
				14'b00010000101110: oled_data = 16'b1111111111111111;
				14'b00010010101110: oled_data = 16'b1111111111111111;
				14'b00010100101110: oled_data = 16'b1111111111111111;
				14'b00010110101110: oled_data = 16'b1111111111111111;
				14'b00011000101110: oled_data = 16'b1111111111111111;
				14'b00011010101110: oled_data = 16'b1111111111111111;
				14'b00011100101110: oled_data = 16'b1111111111111111;
				14'b00011110101110: oled_data = 16'b1111111111111111;
				14'b00100000101110: oled_data = 16'b1111111111111111;
				14'b00100010101110: oled_data = 16'b1111111111111111;
				14'b00100100101110: oled_data = 16'b1111111111111111;
				14'b00100110101110: oled_data = 16'b1111111111111111;
				14'b00101000101110: oled_data = 16'b1111111111111111;
				14'b00101010101110: oled_data = 16'b1111111111111111;
				14'b00101100101110: oled_data = 16'b1111111111111111;
				14'b00101110101110: oled_data = 16'b1111111111111111;
				14'b00110000101110: oled_data = 16'b1111111111111111;
				14'b00110010101110: oled_data = 16'b1111111111111111;
				14'b00110100101110: oled_data = 16'b1111111111111111;
				14'b00110110101110: oled_data = 16'b1111111111111111;
				14'b00111000101110: oled_data = 16'b1111111111111111;
				14'b00111010101110: oled_data = 16'b1111111111111111;
				14'b00111100101110: oled_data = 16'b1111111111111111;
				14'b00111110101110: oled_data = 16'b1111111111111111;
				14'b01000000101110: oled_data = 16'b1111111111111111;
				14'b01000010101110: oled_data = 16'b1111111111111111;
				14'b01000100101110: oled_data = 16'b1111111111111111;
				14'b01000110101110: oled_data = 16'b1111111111111111;
				14'b01001000101110: oled_data = 16'b1111111111111111;
				14'b01001010101110: oled_data = 16'b1111111111111111;
				14'b01001100101110: oled_data = 16'b1111111111111111;
				14'b01001110101110: oled_data = 16'b1111111111111111;
				14'b01010000101110: oled_data = 16'b1111111111111111;
				14'b01010010101110: oled_data = 16'b1111111111111111;
				14'b01010100101110: oled_data = 16'b1111111111111111;
				14'b01010110101110: oled_data = 16'b1111111111111111;
				14'b01011000101110: oled_data = 16'b1111111111111111;
				14'b01011010101110: oled_data = 16'b1111111111111111;
				14'b01011100101110: oled_data = 16'b1111111111111111;
				14'b01011110101110: oled_data = 16'b1111111111111111;
				14'b01100000101110: oled_data = 16'b1111111111111111;
				14'b01100010101110: oled_data = 16'b1111111111111111;
				14'b01100100101110: oled_data = 16'b1111111111111111;
				14'b01100110101110: oled_data = 16'b1111111111111111;
				14'b01101000101110: oled_data = 16'b1111111111111111;
				14'b01101010101110: oled_data = 16'b1111111111111111;
				14'b01101100101110: oled_data = 16'b1111111111111111;
				14'b01101110101110: oled_data = 16'b1111111111111111;
				14'b01110000101110: oled_data = 16'b1111111111111111;
				14'b01110010101110: oled_data = 16'b1111111111111111;
				14'b01110100101110: oled_data = 16'b1111111111111111;
				14'b01110110101110: oled_data = 16'b1111111111111111;
				14'b01111000101110: oled_data = 16'b1111111111111111;
				14'b01111010101110: oled_data = 16'b1111111111111111;
				14'b01111100101110: oled_data = 16'b1111111111111111;
				14'b01111110101110: oled_data = 16'b1111111111111111;
				14'b10000000101110: oled_data = 16'b1111111111111111;
				14'b10000010101110: oled_data = 16'b1111111111111111;
				14'b10000100101110: oled_data = 16'b1111111111111111;
				14'b10000110101110: oled_data = 16'b1111111111111111;
				14'b10001000101110: oled_data = 16'b1111111111111111;
				14'b10001010101110: oled_data = 16'b1111111111111111;
				14'b10001100101110: oled_data = 16'b1111111111111111;
				14'b10001110101110: oled_data = 16'b1111111111111111;
				14'b10010000101110: oled_data = 16'b1111111111111111;
				14'b10010010101110: oled_data = 16'b1111111111111111;
				14'b10010100101110: oled_data = 16'b1111111111111111;
				14'b10010110101110: oled_data = 16'b1111111111111111;
				14'b10011000101110: oled_data = 16'b1111111111111111;
				14'b10011010101110: oled_data = 16'b1111111111111111;
				14'b10011100101110: oled_data = 16'b1111111111111111;
				14'b10011110101110: oled_data = 16'b1111111111111111;
				14'b10100000101110: oled_data = 16'b1111111111111111;
				14'b10100010101110: oled_data = 16'b1111111111111111;
				14'b10100100101110: oled_data = 16'b1111111111111111;
				14'b10100110101110: oled_data = 16'b1111111111111111;
				14'b10101000101110: oled_data = 16'b1111111111111111;
				14'b10101010101110: oled_data = 16'b1111111111111111;
				14'b10101100101110: oled_data = 16'b1111111111111111;
				14'b10101110101110: oled_data = 16'b1111111111111111;
				14'b10110000101110: oled_data = 16'b1111111111111111;
				14'b10110010101110: oled_data = 16'b1111111111111111;
				14'b10110100101110: oled_data = 16'b1111111111111111;
				14'b10110110101110: oled_data = 16'b1111111111111111;
				14'b10111000101110: oled_data = 16'b1111111111111111;
				14'b10111010101110: oled_data = 16'b1111111111111111;
				14'b10111100101110: oled_data = 16'b1111111111111111;
				14'b10111110101110: oled_data = 16'b1111111111111111;
				14'b00000000101111: oled_data = 16'b1111011111011110;
				14'b00000010101111: oled_data = 16'b1110111110111110;
				14'b00000100101111: oled_data = 16'b1110111110011110;
				14'b00000110101111: oled_data = 16'b1110111110011110;
				14'b00001000101111: oled_data = 16'b1110111110011110;
				14'b00001010101111: oled_data = 16'b1110111110111110;
				14'b00001100101111: oled_data = 16'b1110111110111110;
				14'b00001110101111: oled_data = 16'b1111011111011110;
				14'b00010000101111: oled_data = 16'b1111011111011110;
				14'b00010010101111: oled_data = 16'b1111111111111111;
				14'b00010100101111: oled_data = 16'b1111111111111111;
				14'b00010110101111: oled_data = 16'b1111111111111111;
				14'b00011000101111: oled_data = 16'b1111111111111111;
				14'b00011010101111: oled_data = 16'b1111111111111111;
				14'b00011100101111: oled_data = 16'b1111111111111111;
				14'b00011110101111: oled_data = 16'b1111111111111111;
				14'b00100000101111: oled_data = 16'b1111111111111111;
				14'b00100010101111: oled_data = 16'b1111111111111111;
				14'b00100100101111: oled_data = 16'b1111111111111111;
				14'b00100110101111: oled_data = 16'b1111111111111111;
				14'b00101000101111: oled_data = 16'b1111111111111111;
				14'b00101010101111: oled_data = 16'b1111111111111111;
				14'b00101100101111: oled_data = 16'b1111111111111111;
				14'b00101110101111: oled_data = 16'b1111111111111111;
				14'b00110000101111: oled_data = 16'b1111111111111111;
				14'b00110010101111: oled_data = 16'b1111111111111111;
				14'b00110100101111: oled_data = 16'b1111111111111111;
				14'b00110110101111: oled_data = 16'b1111111111111111;
				14'b00111000101111: oled_data = 16'b1111111111111111;
				14'b00111010101111: oled_data = 16'b1111111111111111;
				14'b00111100101111: oled_data = 16'b1111111111111111;
				14'b00111110101111: oled_data = 16'b1111111111111111;
				14'b01000000101111: oled_data = 16'b1111111111111111;
				14'b01000010101111: oled_data = 16'b1111111111111111;
				14'b01000100101111: oled_data = 16'b1111111111111111;
				14'b01000110101111: oled_data = 16'b1111111111111111;
				14'b01001000101111: oled_data = 16'b1111111111111111;
				14'b01001010101111: oled_data = 16'b1111111111111111;
				14'b01001100101111: oled_data = 16'b1111111111111111;
				14'b01001110101111: oled_data = 16'b1111111111111111;
				14'b01010000101111: oled_data = 16'b1111111111111111;
				14'b01010010101111: oled_data = 16'b1111111111111111;
				14'b01010100101111: oled_data = 16'b1111111111111111;
				14'b01010110101111: oled_data = 16'b1111111111111111;
				14'b01011000101111: oled_data = 16'b1111111111111111;
				14'b01011010101111: oled_data = 16'b1111111111111111;
				14'b01011100101111: oled_data = 16'b1111111111111111;
				14'b01011110101111: oled_data = 16'b1111111111111111;
				14'b01100000101111: oled_data = 16'b1111111111111111;
				14'b01100010101111: oled_data = 16'b1111111111111111;
				14'b01100100101111: oled_data = 16'b1111111111111111;
				14'b01100110101111: oled_data = 16'b1111111111111111;
				14'b01101000101111: oled_data = 16'b1111111111111111;
				14'b01101010101111: oled_data = 16'b1111111111111111;
				14'b01101100101111: oled_data = 16'b1111111111111111;
				14'b01101110101111: oled_data = 16'b1111111111111111;
				14'b01110000101111: oled_data = 16'b1111111111111111;
				14'b01110010101111: oled_data = 16'b1111111111111111;
				14'b01110100101111: oled_data = 16'b1111111111111111;
				14'b01110110101111: oled_data = 16'b1111111111111111;
				14'b01111000101111: oled_data = 16'b1111111111111111;
				14'b01111010101111: oled_data = 16'b1111111111111111;
				14'b01111100101111: oled_data = 16'b1111111111111111;
				14'b01111110101111: oled_data = 16'b1111111111111111;
				14'b10000000101111: oled_data = 16'b1111111111111111;
				14'b10000010101111: oled_data = 16'b1111111111111111;
				14'b10000100101111: oled_data = 16'b1111111111111111;
				14'b10000110101111: oled_data = 16'b1111111111111111;
				14'b10001000101111: oled_data = 16'b1111111111111111;
				14'b10001010101111: oled_data = 16'b1111111111111111;
				14'b10001100101111: oled_data = 16'b1111111111111111;
				14'b10001110101111: oled_data = 16'b1111111111111111;
				14'b10010000101111: oled_data = 16'b1111111111111111;
				14'b10010010101111: oled_data = 16'b1111111111111111;
				14'b10010100101111: oled_data = 16'b1111111111111111;
				14'b10010110101111: oled_data = 16'b1111111111111111;
				14'b10011000101111: oled_data = 16'b1111111111111111;
				14'b10011010101111: oled_data = 16'b1111111111111111;
				14'b10011100101111: oled_data = 16'b1111111111111111;
				14'b10011110101111: oled_data = 16'b1111111111111111;
				14'b10100000101111: oled_data = 16'b1111111111111111;
				14'b10100010101111: oled_data = 16'b1111111111111111;
				14'b10100100101111: oled_data = 16'b1111111111111111;
				14'b10100110101111: oled_data = 16'b1111111111111111;
				14'b10101000101111: oled_data = 16'b1111111111111111;
				14'b10101010101111: oled_data = 16'b1111111111111111;
				14'b10101100101111: oled_data = 16'b1111111111111111;
				14'b10101110101111: oled_data = 16'b1111111111111111;
				14'b10110000101111: oled_data = 16'b1111111111111111;
				14'b10110010101111: oled_data = 16'b1111111111111111;
				14'b10110100101111: oled_data = 16'b1111111111111111;
				14'b10110110101111: oled_data = 16'b1111111111111111;
				14'b10111000101111: oled_data = 16'b1111111111111111;
				14'b10111010101111: oled_data = 16'b1111111111111111;
				14'b10111100101111: oled_data = 16'b1111111111111111;
				14'b10111110101111: oled_data = 16'b1111111111111111;
				14'b00000000110000: oled_data = 16'b1101111100111101;
				14'b00000010110000: oled_data = 16'b1101011100011100;
				14'b00000100110000: oled_data = 16'b1101011100011100;
				14'b00000110110000: oled_data = 16'b1101011100011100;
				14'b00001000110000: oled_data = 16'b1101011100011100;
				14'b00001010110000: oled_data = 16'b1101111100111100;
				14'b00001100110000: oled_data = 16'b1101111101011100;
				14'b00001110110000: oled_data = 16'b1110011110011101;
				14'b00010000110000: oled_data = 16'b1110111110111101;
				14'b00010010110000: oled_data = 16'b1111011111011110;
				14'b00010100110000: oled_data = 16'b1111011111011110;
				14'b00010110110000: oled_data = 16'b1111111111111111;
				14'b00011000110000: oled_data = 16'b1111111111111111;
				14'b00011010110000: oled_data = 16'b1111111111111111;
				14'b00011100110000: oled_data = 16'b1111111111111111;
				14'b00011110110000: oled_data = 16'b1111111111111111;
				14'b00100000110000: oled_data = 16'b1111111111111111;
				14'b00100010110000: oled_data = 16'b1111111111111111;
				14'b00100100110000: oled_data = 16'b1111111111111111;
				14'b00100110110000: oled_data = 16'b1111111111111111;
				14'b00101000110000: oled_data = 16'b1111111111111111;
				14'b00101010110000: oled_data = 16'b1111111111111111;
				14'b00101100110000: oled_data = 16'b1111111111111111;
				14'b00101110110000: oled_data = 16'b1111111111111111;
				14'b00110000110000: oled_data = 16'b1111111111111111;
				14'b00110010110000: oled_data = 16'b1111111111111111;
				14'b00110100110000: oled_data = 16'b1111111111111111;
				14'b00110110110000: oled_data = 16'b1111111111111111;
				14'b00111000110000: oled_data = 16'b1111111111111111;
				14'b00111010110000: oled_data = 16'b1111111111111111;
				14'b00111100110000: oled_data = 16'b1111111111111111;
				14'b00111110110000: oled_data = 16'b1111111111111111;
				14'b01000000110000: oled_data = 16'b1111111111111111;
				14'b01000010110000: oled_data = 16'b1111111111111111;
				14'b01000100110000: oled_data = 16'b1111111111111111;
				14'b01000110110000: oled_data = 16'b1111111111111111;
				14'b01001000110000: oled_data = 16'b1111111111111111;
				14'b01001010110000: oled_data = 16'b1111111111111111;
				14'b01001100110000: oled_data = 16'b1111111111111111;
				14'b01001110110000: oled_data = 16'b1111111111111111;
				14'b01010000110000: oled_data = 16'b1111111111111111;
				14'b01010010110000: oled_data = 16'b1111111111111111;
				14'b01010100110000: oled_data = 16'b1111111111111111;
				14'b01010110110000: oled_data = 16'b1111111111111111;
				14'b01011000110000: oled_data = 16'b1111111111111111;
				14'b01011010110000: oled_data = 16'b1111111111111111;
				14'b01011100110000: oled_data = 16'b1111111111111111;
				14'b01011110110000: oled_data = 16'b1111111111111111;
				14'b01100000110000: oled_data = 16'b1111111111111111;
				14'b01100010110000: oled_data = 16'b1111111111111111;
				14'b01100100110000: oled_data = 16'b1111111111111111;
				14'b01100110110000: oled_data = 16'b1111111111111111;
				14'b01101000110000: oled_data = 16'b1111111111111111;
				14'b01101010110000: oled_data = 16'b1111111111111111;
				14'b01101100110000: oled_data = 16'b1111111111111111;
				14'b01101110110000: oled_data = 16'b1111111111111111;
				14'b01110000110000: oled_data = 16'b1111111111111111;
				14'b01110010110000: oled_data = 16'b1111111111111111;
				14'b01110100110000: oled_data = 16'b1111111111111111;
				14'b01110110110000: oled_data = 16'b1111111111111111;
				14'b01111000110000: oled_data = 16'b1111111111111111;
				14'b01111010110000: oled_data = 16'b1111111111111111;
				14'b01111100110000: oled_data = 16'b1111111111111111;
				14'b01111110110000: oled_data = 16'b1111111111111111;
				14'b10000000110000: oled_data = 16'b1111111111111111;
				14'b10000010110000: oled_data = 16'b1111111111111111;
				14'b10000100110000: oled_data = 16'b1111111111111111;
				14'b10000110110000: oled_data = 16'b1111111111111111;
				14'b10001000110000: oled_data = 16'b1111111111111111;
				14'b10001010110000: oled_data = 16'b1111111111111111;
				14'b10001100110000: oled_data = 16'b1111111111111111;
				14'b10001110110000: oled_data = 16'b1111111111111111;
				14'b10010000110000: oled_data = 16'b1111111111111111;
				14'b10010010110000: oled_data = 16'b1111111111111111;
				14'b10010100110000: oled_data = 16'b1111111111111111;
				14'b10010110110000: oled_data = 16'b1111111111111111;
				14'b10011000110000: oled_data = 16'b1111111111111111;
				14'b10011010110000: oled_data = 16'b1111111111111111;
				14'b10011100110000: oled_data = 16'b1111111111111111;
				14'b10011110110000: oled_data = 16'b1111111111111111;
				14'b10100000110000: oled_data = 16'b1111111111111111;
				14'b10100010110000: oled_data = 16'b1111111111111111;
				14'b10100100110000: oled_data = 16'b1111111111111111;
				14'b10100110110000: oled_data = 16'b1111111111111111;
				14'b10101000110000: oled_data = 16'b1111111111111111;
				14'b10101010110000: oled_data = 16'b1111111111111111;
				14'b10101100110000: oled_data = 16'b1111111111111111;
				14'b10101110110000: oled_data = 16'b1111111111111111;
				14'b10110000110000: oled_data = 16'b1111111111111111;
				14'b10110010110000: oled_data = 16'b1111111111111111;
				14'b10110100110000: oled_data = 16'b1111111111111111;
				14'b10110110110000: oled_data = 16'b1111111111111111;
				14'b10111000110000: oled_data = 16'b1111111111111111;
				14'b10111010110000: oled_data = 16'b1111111111111111;
				14'b10111100110000: oled_data = 16'b1111111111111111;
				14'b10111110110000: oled_data = 16'b1111111111111111;
				14'b00000000110001: oled_data = 16'b1100011010111100;
				14'b00000010110001: oled_data = 16'b1100111011011100;
				14'b00000100110001: oled_data = 16'b1100111011011100;
				14'b00000110110001: oled_data = 16'b1100111011011011;
				14'b00001000110001: oled_data = 16'b1100111011111011;
				14'b00001010110001: oled_data = 16'b1100111011011011;
				14'b00001100110001: oled_data = 16'b1100111011011010;
				14'b00001110110001: oled_data = 16'b1100111100011011;
				14'b00010000110001: oled_data = 16'b1101011100111011;
				14'b00010010110001: oled_data = 16'b1110011101111100;
				14'b00010100110001: oled_data = 16'b1110111110111101;
				14'b00010110110001: oled_data = 16'b1111011111011110;
				14'b00011000110001: oled_data = 16'b1111111111111111;
				14'b00011010110001: oled_data = 16'b1111111111111111;
				14'b00011100110001: oled_data = 16'b1111111111111111;
				14'b00011110110001: oled_data = 16'b1111111111111111;
				14'b00100000110001: oled_data = 16'b1111111111111111;
				14'b00100010110001: oled_data = 16'b1111111111111111;
				14'b00100100110001: oled_data = 16'b1111111111111111;
				14'b00100110110001: oled_data = 16'b1111111111111111;
				14'b00101000110001: oled_data = 16'b1111111111111111;
				14'b00101010110001: oled_data = 16'b1111111111111111;
				14'b00101100110001: oled_data = 16'b1111111111111111;
				14'b00101110110001: oled_data = 16'b1111111111111111;
				14'b00110000110001: oled_data = 16'b1111111111111111;
				14'b00110010110001: oled_data = 16'b1111111111111111;
				14'b00110100110001: oled_data = 16'b1111111111111111;
				14'b00110110110001: oled_data = 16'b1111111111111111;
				14'b00111000110001: oled_data = 16'b1111111111111111;
				14'b00111010110001: oled_data = 16'b1111111111111111;
				14'b00111100110001: oled_data = 16'b1111111111111111;
				14'b00111110110001: oled_data = 16'b1111111111111111;
				14'b01000000110001: oled_data = 16'b1111111111111111;
				14'b01000010110001: oled_data = 16'b1111111111111111;
				14'b01000100110001: oled_data = 16'b1111111111111111;
				14'b01000110110001: oled_data = 16'b1111111111111111;
				14'b01001000110001: oled_data = 16'b1111111111111111;
				14'b01001010110001: oled_data = 16'b1111111111111111;
				14'b01001100110001: oled_data = 16'b1111111111111111;
				14'b01001110110001: oled_data = 16'b1111111111111111;
				14'b01010000110001: oled_data = 16'b1111111111111111;
				14'b01010010110001: oled_data = 16'b1111111111111111;
				14'b01010100110001: oled_data = 16'b1111111111111111;
				14'b01010110110001: oled_data = 16'b1111111111111111;
				14'b01011000110001: oled_data = 16'b1111111111111111;
				14'b01011010110001: oled_data = 16'b1111111111111111;
				14'b01011100110001: oled_data = 16'b1111111111111111;
				14'b01011110110001: oled_data = 16'b1111111111111111;
				14'b01100000110001: oled_data = 16'b1111111111111111;
				14'b01100010110001: oled_data = 16'b1111111111111111;
				14'b01100100110001: oled_data = 16'b1111111111111111;
				14'b01100110110001: oled_data = 16'b1111111111111111;
				14'b01101000110001: oled_data = 16'b1111111111111111;
				14'b01101010110001: oled_data = 16'b1111111111111111;
				14'b01101100110001: oled_data = 16'b1111111111111111;
				14'b01101110110001: oled_data = 16'b1111111111111111;
				14'b01110000110001: oled_data = 16'b1111111111111111;
				14'b01110010110001: oled_data = 16'b1111111111111111;
				14'b01110100110001: oled_data = 16'b1111111111111111;
				14'b01110110110001: oled_data = 16'b1111111111111111;
				14'b01111000110001: oled_data = 16'b1111111111111111;
				14'b01111010110001: oled_data = 16'b1111111111111111;
				14'b01111100110001: oled_data = 16'b1111111111111111;
				14'b01111110110001: oled_data = 16'b1111111111111111;
				14'b10000000110001: oled_data = 16'b1111111111111111;
				14'b10000010110001: oled_data = 16'b1111111111111111;
				14'b10000100110001: oled_data = 16'b1111111111111111;
				14'b10000110110001: oled_data = 16'b1111111111111111;
				14'b10001000110001: oled_data = 16'b1111111111111111;
				14'b10001010110001: oled_data = 16'b1111111111111111;
				14'b10001100110001: oled_data = 16'b1111111111111111;
				14'b10001110110001: oled_data = 16'b1111111111111111;
				14'b10010000110001: oled_data = 16'b1111111111111111;
				14'b10010010110001: oled_data = 16'b1111111111111111;
				14'b10010100110001: oled_data = 16'b1111111111111111;
				14'b10010110110001: oled_data = 16'b1111111111111111;
				14'b10011000110001: oled_data = 16'b1111111111111111;
				14'b10011010110001: oled_data = 16'b1111111111111111;
				14'b10011100110001: oled_data = 16'b1111111111111111;
				14'b10011110110001: oled_data = 16'b1111111111111111;
				14'b10100000110001: oled_data = 16'b1111111111111111;
				14'b10100010110001: oled_data = 16'b1111111111111111;
				14'b10100100110001: oled_data = 16'b1111111111111111;
				14'b10100110110001: oled_data = 16'b1111111111111111;
				14'b10101000110001: oled_data = 16'b1111111111111111;
				14'b10101010110001: oled_data = 16'b1111111111111111;
				14'b10101100110001: oled_data = 16'b1111111111111111;
				14'b10101110110001: oled_data = 16'b1111111111111111;
				14'b10110000110001: oled_data = 16'b1111111111111111;
				14'b10110010110001: oled_data = 16'b1111111111111111;
				14'b10110100110001: oled_data = 16'b1111111111111111;
				14'b10110110110001: oled_data = 16'b1111111111111111;
				14'b10111000110001: oled_data = 16'b1111111111111111;
				14'b10111010110001: oled_data = 16'b1111111111111111;
				14'b10111100110001: oled_data = 16'b1111111111111111;
				14'b10111110110001: oled_data = 16'b1111111111111111;
				14'b00000000110010: oled_data = 16'b1101011011111101;
				14'b00000010110010: oled_data = 16'b1101011100011101;
				14'b00000100110010: oled_data = 16'b1101011100011100;
				14'b00000110110010: oled_data = 16'b1101011100011100;
				14'b00001000110010: oled_data = 16'b1101011100111100;
				14'b00001010110010: oled_data = 16'b1101011100111100;
				14'b00001100110010: oled_data = 16'b1101011100011011;
				14'b00001110110010: oled_data = 16'b1101011100011011;
				14'b00010000110010: oled_data = 16'b1100111100011010;
				14'b00010010110010: oled_data = 16'b1100111100011010;
				14'b00010100110010: oled_data = 16'b1101011100111011;
				14'b00010110110010: oled_data = 16'b1110011110011100;
				14'b00011000110010: oled_data = 16'b1111011111011110;
				14'b00011010110010: oled_data = 16'b1111111111111111;
				14'b00011100110010: oled_data = 16'b1111111111111111;
				14'b00011110110010: oled_data = 16'b1111111111111111;
				14'b00100000110010: oled_data = 16'b1111111111111111;
				14'b00100010110010: oled_data = 16'b1111111111111111;
				14'b00100100110010: oled_data = 16'b1111111111111111;
				14'b00100110110010: oled_data = 16'b1111111111111111;
				14'b00101000110010: oled_data = 16'b1111111111111111;
				14'b00101010110010: oled_data = 16'b1111111111111111;
				14'b00101100110010: oled_data = 16'b1111111111111111;
				14'b00101110110010: oled_data = 16'b1111111111111111;
				14'b00110000110010: oled_data = 16'b1111111111111111;
				14'b00110010110010: oled_data = 16'b1111111111111111;
				14'b00110100110010: oled_data = 16'b1111111111111111;
				14'b00110110110010: oled_data = 16'b1111111111111111;
				14'b00111000110010: oled_data = 16'b1111111111111111;
				14'b00111010110010: oled_data = 16'b1111111111111111;
				14'b00111100110010: oled_data = 16'b1111111111111111;
				14'b00111110110010: oled_data = 16'b1111111111111111;
				14'b01000000110010: oled_data = 16'b1111111111111111;
				14'b01000010110010: oled_data = 16'b1111111111111111;
				14'b01000100110010: oled_data = 16'b1111111111111111;
				14'b01000110110010: oled_data = 16'b1111111111111111;
				14'b01001000110010: oled_data = 16'b1111111111111111;
				14'b01001010110010: oled_data = 16'b1111111111111111;
				14'b01001100110010: oled_data = 16'b1111111111111111;
				14'b01001110110010: oled_data = 16'b1111111111111111;
				14'b01010000110010: oled_data = 16'b1111111111111111;
				14'b01010010110010: oled_data = 16'b1111111111111111;
				14'b01010100110010: oled_data = 16'b1111111111111111;
				14'b01010110110010: oled_data = 16'b1111111111111111;
				14'b01011000110010: oled_data = 16'b1111111111111111;
				14'b01011010110010: oled_data = 16'b1111111111111111;
				14'b01011100110010: oled_data = 16'b1111111111111111;
				14'b01011110110010: oled_data = 16'b1111111111111111;
				14'b01100000110010: oled_data = 16'b1111111111111111;
				14'b01100010110010: oled_data = 16'b1111111111111111;
				14'b01100100110010: oled_data = 16'b1111111111111111;
				14'b01100110110010: oled_data = 16'b1111111111111111;
				14'b01101000110010: oled_data = 16'b1111111111111111;
				14'b01101010110010: oled_data = 16'b1111111111111111;
				14'b01101100110010: oled_data = 16'b1111111111111111;
				14'b01101110110010: oled_data = 16'b1111111111111111;
				14'b01110000110010: oled_data = 16'b1111111111111111;
				14'b01110010110010: oled_data = 16'b1111111111111111;
				14'b01110100110010: oled_data = 16'b1111111111111111;
				14'b01110110110010: oled_data = 16'b1111111111111111;
				14'b01111000110010: oled_data = 16'b1111111111111111;
				14'b01111010110010: oled_data = 16'b1111111111111111;
				14'b01111100110010: oled_data = 16'b1111111111111111;
				14'b01111110110010: oled_data = 16'b1111111111111111;
				14'b10000000110010: oled_data = 16'b1111111111111111;
				14'b10000010110010: oled_data = 16'b1111111111111111;
				14'b10000100110010: oled_data = 16'b1111111111111111;
				14'b10000110110010: oled_data = 16'b1111111111111111;
				14'b10001000110010: oled_data = 16'b1111111111111111;
				14'b10001010110010: oled_data = 16'b1111111111111111;
				14'b10001100110010: oled_data = 16'b1111111111111111;
				14'b10001110110010: oled_data = 16'b1111111111111111;
				14'b10010000110010: oled_data = 16'b1111111111111111;
				14'b10010010110010: oled_data = 16'b1111111111111111;
				14'b10010100110010: oled_data = 16'b1111111111111111;
				14'b10010110110010: oled_data = 16'b1111111111111111;
				14'b10011000110010: oled_data = 16'b1111111111111111;
				14'b10011010110010: oled_data = 16'b1111111111111111;
				14'b10011100110010: oled_data = 16'b1111111111111111;
				14'b10011110110010: oled_data = 16'b1111111111111111;
				14'b10100000110010: oled_data = 16'b1111111111111111;
				14'b10100010110010: oled_data = 16'b1111111111111111;
				14'b10100100110010: oled_data = 16'b1111111111111111;
				14'b10100110110010: oled_data = 16'b1111111111111111;
				14'b10101000110010: oled_data = 16'b1111111111111111;
				14'b10101010110010: oled_data = 16'b1111111111111111;
				14'b10101100110010: oled_data = 16'b1111111111111111;
				14'b10101110110010: oled_data = 16'b1111111111111111;
				14'b10110000110010: oled_data = 16'b1111111111111111;
				14'b10110010110010: oled_data = 16'b1111111111111111;
				14'b10110100110010: oled_data = 16'b1111111111111111;
				14'b10110110110010: oled_data = 16'b1111111111111111;
				14'b10111000110010: oled_data = 16'b1111111111111111;
				14'b10111010110010: oled_data = 16'b1111111111111111;
				14'b10111100110010: oled_data = 16'b1111111111111111;
				14'b10111110110010: oled_data = 16'b1111111111111111;
				14'b00000000110011: oled_data = 16'b1101111101011101;
				14'b00000010110011: oled_data = 16'b1110011101111101;
				14'b00000100110011: oled_data = 16'b1110011101111101;
				14'b00000110110011: oled_data = 16'b1110011101111101;
				14'b00001000110011: oled_data = 16'b1110011101111101;
				14'b00001010110011: oled_data = 16'b1101111101011101;
				14'b00001100110011: oled_data = 16'b1101111100111100;
				14'b00001110110011: oled_data = 16'b1101111100111100;
				14'b00010000110011: oled_data = 16'b1101111100111100;
				14'b00010010110011: oled_data = 16'b1101011100111011;
				14'b00010100110011: oled_data = 16'b1100111100011010;
				14'b00010110110011: oled_data = 16'b1101011100011010;
				14'b00011000110011: oled_data = 16'b1101111101111011;
				14'b00011010110011: oled_data = 16'b1111011110111110;
				14'b00011100110011: oled_data = 16'b1111111111111111;
				14'b00011110110011: oled_data = 16'b1111111111111111;
				14'b00100000110011: oled_data = 16'b1111111111111111;
				14'b00100010110011: oled_data = 16'b1111111111111111;
				14'b00100100110011: oled_data = 16'b1111111111111111;
				14'b00100110110011: oled_data = 16'b1111111111111111;
				14'b00101000110011: oled_data = 16'b1111111111111111;
				14'b00101010110011: oled_data = 16'b1111111111111111;
				14'b00101100110011: oled_data = 16'b1111111111111111;
				14'b00101110110011: oled_data = 16'b1111111111111111;
				14'b00110000110011: oled_data = 16'b1111111111111111;
				14'b00110010110011: oled_data = 16'b1111111111111111;
				14'b00110100110011: oled_data = 16'b1111111111111111;
				14'b00110110110011: oled_data = 16'b1111111111111111;
				14'b00111000110011: oled_data = 16'b1111111111111111;
				14'b00111010110011: oled_data = 16'b1111111111111111;
				14'b00111100110011: oled_data = 16'b1111111111111111;
				14'b00111110110011: oled_data = 16'b1111111111111111;
				14'b01000000110011: oled_data = 16'b1111111111111111;
				14'b01000010110011: oled_data = 16'b1111111111111111;
				14'b01000100110011: oled_data = 16'b1111111111111111;
				14'b01000110110011: oled_data = 16'b1111111111111111;
				14'b01001000110011: oled_data = 16'b1111111111111111;
				14'b01001010110011: oled_data = 16'b1111111111111111;
				14'b01001100110011: oled_data = 16'b1111111111111111;
				14'b01001110110011: oled_data = 16'b1111111111111111;
				14'b01010000110011: oled_data = 16'b1111111111111111;
				14'b01010010110011: oled_data = 16'b1111111111111111;
				14'b01010100110011: oled_data = 16'b1111111111111111;
				14'b01010110110011: oled_data = 16'b1111111111111111;
				14'b01011000110011: oled_data = 16'b1111111111111111;
				14'b01011010110011: oled_data = 16'b1111111111111111;
				14'b01011100110011: oled_data = 16'b1111111111111111;
				14'b01011110110011: oled_data = 16'b1111111111111111;
				14'b01100000110011: oled_data = 16'b1111111111111111;
				14'b01100010110011: oled_data = 16'b1111111111111111;
				14'b01100100110011: oled_data = 16'b1111111111111111;
				14'b01100110110011: oled_data = 16'b1111111111111111;
				14'b01101000110011: oled_data = 16'b1111111111111111;
				14'b01101010110011: oled_data = 16'b1111111111111111;
				14'b01101100110011: oled_data = 16'b1111111111111111;
				14'b01101110110011: oled_data = 16'b1111111111111111;
				14'b01110000110011: oled_data = 16'b1111111111111111;
				14'b01110010110011: oled_data = 16'b1111111111111111;
				14'b01110100110011: oled_data = 16'b1111111111111111;
				14'b01110110110011: oled_data = 16'b1111111111111111;
				14'b01111000110011: oled_data = 16'b1111111111111111;
				14'b01111010110011: oled_data = 16'b1111111111111111;
				14'b01111100110011: oled_data = 16'b1111111111111111;
				14'b01111110110011: oled_data = 16'b1111111111111111;
				14'b10000000110011: oled_data = 16'b1111111111111111;
				14'b10000010110011: oled_data = 16'b1111111111111111;
				14'b10000100110011: oled_data = 16'b1111111111111111;
				14'b10000110110011: oled_data = 16'b1111111111111111;
				14'b10001000110011: oled_data = 16'b1111111111111111;
				14'b10001010110011: oled_data = 16'b1111111111111111;
				14'b10001100110011: oled_data = 16'b1111111111111111;
				14'b10001110110011: oled_data = 16'b1111111111111111;
				14'b10010000110011: oled_data = 16'b1111111111111111;
				14'b10010010110011: oled_data = 16'b1111111111111111;
				14'b10010100110011: oled_data = 16'b1111111111111111;
				14'b10010110110011: oled_data = 16'b1111111111111111;
				14'b10011000110011: oled_data = 16'b1111111111111111;
				14'b10011010110011: oled_data = 16'b1111111111111111;
				14'b10011100110011: oled_data = 16'b1111111111111111;
				14'b10011110110011: oled_data = 16'b1111111111111111;
				14'b10100000110011: oled_data = 16'b1111111111111111;
				14'b10100010110011: oled_data = 16'b1111111111111111;
				14'b10100100110011: oled_data = 16'b1111111111111111;
				14'b10100110110011: oled_data = 16'b1111111111111111;
				14'b10101000110011: oled_data = 16'b1111111111111111;
				14'b10101010110011: oled_data = 16'b1111111111111111;
				14'b10101100110011: oled_data = 16'b1111111111111111;
				14'b10101110110011: oled_data = 16'b1111111111111111;
				14'b10110000110011: oled_data = 16'b1111111111111111;
				14'b10110010110011: oled_data = 16'b1111111111111111;
				14'b10110100110011: oled_data = 16'b1111111111111111;
				14'b10110110110011: oled_data = 16'b1111111111111111;
				14'b10111000110011: oled_data = 16'b1111111111111111;
				14'b10111010110011: oled_data = 16'b1111111111111111;
				14'b10111100110011: oled_data = 16'b1111111111111111;
				14'b10111110110011: oled_data = 16'b1111111111111111;
				14'b00000000110100: oled_data = 16'b1111011111011110;
				14'b00000010110100: oled_data = 16'b1111111111111111;
				14'b00000100110100: oled_data = 16'b1111111111111111;
				14'b00000110110100: oled_data = 16'b1111111111111111;
				14'b00001000110100: oled_data = 16'b1111111111111111;
				14'b00001010110100: oled_data = 16'b1111011111011110;
				14'b00001100110100: oled_data = 16'b1111011110111110;
				14'b00001110110100: oled_data = 16'b1110111110011101;
				14'b00010000110100: oled_data = 16'b1101111101011100;
				14'b00010010110100: oled_data = 16'b1101111101011100;
				14'b00010100110100: oled_data = 16'b1101111101011011;
				14'b00010110110100: oled_data = 16'b1101011100111010;
				14'b00011000110100: oled_data = 16'b1100111100011001;
				14'b00011010110100: oled_data = 16'b1101111101011011;
				14'b00011100110100: oled_data = 16'b1111011111011110;
				14'b00011110110100: oled_data = 16'b1111111111111111;
				14'b00100000110100: oled_data = 16'b1111111111111111;
				14'b00100010110100: oled_data = 16'b1111111111111111;
				14'b00100100110100: oled_data = 16'b1111111111111111;
				14'b00100110110100: oled_data = 16'b1111111111111111;
				14'b00101000110100: oled_data = 16'b1111111111111111;
				14'b00101010110100: oled_data = 16'b1111111111111111;
				14'b00101100110100: oled_data = 16'b1111111111111111;
				14'b00101110110100: oled_data = 16'b1111111111111111;
				14'b00110000110100: oled_data = 16'b1111111111111111;
				14'b00110010110100: oled_data = 16'b1111111111111111;
				14'b00110100110100: oled_data = 16'b1111111111111111;
				14'b00110110110100: oled_data = 16'b1111111111111111;
				14'b00111000110100: oled_data = 16'b1111111111111111;
				14'b00111010110100: oled_data = 16'b1111111111111111;
				14'b00111100110100: oled_data = 16'b1111111111111111;
				14'b00111110110100: oled_data = 16'b1111111111111111;
				14'b01000000110100: oled_data = 16'b1111111111111111;
				14'b01000010110100: oled_data = 16'b1111111111111111;
				14'b01000100110100: oled_data = 16'b1111111111111111;
				14'b01000110110100: oled_data = 16'b1111111111111111;
				14'b01001000110100: oled_data = 16'b1111111111111111;
				14'b01001010110100: oled_data = 16'b1111111111111111;
				14'b01001100110100: oled_data = 16'b1111111111111111;
				14'b01001110110100: oled_data = 16'b1111111111111111;
				14'b01010000110100: oled_data = 16'b1111111111111111;
				14'b01010010110100: oled_data = 16'b1111111111111111;
				14'b01010100110100: oled_data = 16'b1111111111111111;
				14'b01010110110100: oled_data = 16'b1111111111111111;
				14'b01011000110100: oled_data = 16'b1111111111111111;
				14'b01011010110100: oled_data = 16'b1111111111111111;
				14'b01011100110100: oled_data = 16'b1111111111111111;
				14'b01011110110100: oled_data = 16'b1111111111111111;
				14'b01100000110100: oled_data = 16'b1111111111111111;
				14'b01100010110100: oled_data = 16'b1111111111111111;
				14'b01100100110100: oled_data = 16'b1111111111111111;
				14'b01100110110100: oled_data = 16'b1111111111111111;
				14'b01101000110100: oled_data = 16'b1111111111111111;
				14'b01101010110100: oled_data = 16'b1111111111111111;
				14'b01101100110100: oled_data = 16'b1111111111111111;
				14'b01101110110100: oled_data = 16'b1111111111111111;
				14'b01110000110100: oled_data = 16'b1111111111111111;
				14'b01110010110100: oled_data = 16'b1111111111111111;
				14'b01110100110100: oled_data = 16'b1111111111111111;
				14'b01110110110100: oled_data = 16'b1111111111111111;
				14'b01111000110100: oled_data = 16'b1111111111111111;
				14'b01111010110100: oled_data = 16'b1111111111111111;
				14'b01111100110100: oled_data = 16'b1111111111111111;
				14'b01111110110100: oled_data = 16'b1111111111111111;
				14'b10000000110100: oled_data = 16'b1111111111111111;
				14'b10000010110100: oled_data = 16'b1111111111111111;
				14'b10000100110100: oled_data = 16'b1111111111111111;
				14'b10000110110100: oled_data = 16'b1111111111111111;
				14'b10001000110100: oled_data = 16'b1111111111111111;
				14'b10001010110100: oled_data = 16'b1111111111111111;
				14'b10001100110100: oled_data = 16'b1111111111111111;
				14'b10001110110100: oled_data = 16'b1111111111111111;
				14'b10010000110100: oled_data = 16'b1111111111111111;
				14'b10010010110100: oled_data = 16'b1111111111111111;
				14'b10010100110100: oled_data = 16'b1111111111111111;
				14'b10010110110100: oled_data = 16'b1111111111111111;
				14'b10011000110100: oled_data = 16'b1111111111111111;
				14'b10011010110100: oled_data = 16'b1111111111111111;
				14'b10011100110100: oled_data = 16'b1111111111111111;
				14'b10011110110100: oled_data = 16'b1111111111111111;
				14'b10100000110100: oled_data = 16'b1111111111111111;
				14'b10100010110100: oled_data = 16'b1111111111111111;
				14'b10100100110100: oled_data = 16'b1111111111111111;
				14'b10100110110100: oled_data = 16'b1111111111111111;
				14'b10101000110100: oled_data = 16'b1111111111111111;
				14'b10101010110100: oled_data = 16'b1111111111111111;
				14'b10101100110100: oled_data = 16'b1111111111111111;
				14'b10101110110100: oled_data = 16'b1111111111111111;
				14'b10110000110100: oled_data = 16'b1111111111111111;
				14'b10110010110100: oled_data = 16'b1111111111111111;
				14'b10110100110100: oled_data = 16'b1111111111111111;
				14'b10110110110100: oled_data = 16'b1111111111111111;
				14'b10111000110100: oled_data = 16'b1111111111111111;
				14'b10111010110100: oled_data = 16'b1111111111111111;
				14'b10111100110100: oled_data = 16'b1111111111111111;
				14'b10111110110100: oled_data = 16'b1111111111111111;
				14'b00000000110101: oled_data = 16'b1111111111111111;
				14'b00000010110101: oled_data = 16'b1111111111111111;
				14'b00000100110101: oled_data = 16'b1111111111111111;
				14'b00000110110101: oled_data = 16'b1111111111111111;
				14'b00001000110101: oled_data = 16'b1111111111111111;
				14'b00001010110101: oled_data = 16'b1111111111111111;
				14'b00001100110101: oled_data = 16'b1111111111111111;
				14'b00001110110101: oled_data = 16'b1111111111111111;
				14'b00010000110101: oled_data = 16'b1111011111011110;
				14'b00010010110101: oled_data = 16'b1110111110011101;
				14'b00010100110101: oled_data = 16'b1101111101011100;
				14'b00010110110101: oled_data = 16'b1101111101011011;
				14'b00011000110101: oled_data = 16'b1101011101011010;
				14'b00011010110101: oled_data = 16'b1100111100011001;
				14'b00011100110101: oled_data = 16'b1101111101011010;
				14'b00011110110101: oled_data = 16'b1111011111011110;
				14'b00100000110101: oled_data = 16'b1111111111111111;
				14'b00100010110101: oled_data = 16'b1111111111111111;
				14'b00100100110101: oled_data = 16'b1111111111111111;
				14'b00100110110101: oled_data = 16'b1111111111111111;
				14'b00101000110101: oled_data = 16'b1111111111111111;
				14'b00101010110101: oled_data = 16'b1111111111111111;
				14'b00101100110101: oled_data = 16'b1111111111111111;
				14'b00101110110101: oled_data = 16'b1111111111111111;
				14'b00110000110101: oled_data = 16'b1111111111111111;
				14'b00110010110101: oled_data = 16'b1111111111111111;
				14'b00110100110101: oled_data = 16'b1111111111111111;
				14'b00110110110101: oled_data = 16'b1111111111111111;
				14'b00111000110101: oled_data = 16'b1111111111111111;
				14'b00111010110101: oled_data = 16'b1111111111111111;
				14'b00111100110101: oled_data = 16'b1111111111111111;
				14'b00111110110101: oled_data = 16'b1111111111111111;
				14'b01000000110101: oled_data = 16'b1111111111111111;
				14'b01000010110101: oled_data = 16'b1111111111111111;
				14'b01000100110101: oled_data = 16'b1111111111111111;
				14'b01000110110101: oled_data = 16'b1111111111111111;
				14'b01001000110101: oled_data = 16'b1111111111111111;
				14'b01001010110101: oled_data = 16'b1111111111111111;
				14'b01001100110101: oled_data = 16'b1111111111111111;
				14'b01001110110101: oled_data = 16'b1111111111111111;
				14'b01010000110101: oled_data = 16'b1111111111111111;
				14'b01010010110101: oled_data = 16'b1111111111111111;
				14'b01010100110101: oled_data = 16'b1111111111111111;
				14'b01010110110101: oled_data = 16'b1111111111111111;
				14'b01011000110101: oled_data = 16'b1111111111111111;
				14'b01011010110101: oled_data = 16'b1111111111111111;
				14'b01011100110101: oled_data = 16'b1111111111111111;
				14'b01011110110101: oled_data = 16'b1111111111111111;
				14'b01100000110101: oled_data = 16'b1111111111111111;
				14'b01100010110101: oled_data = 16'b1111111111111111;
				14'b01100100110101: oled_data = 16'b1111111111111111;
				14'b01100110110101: oled_data = 16'b1111111111111111;
				14'b01101000110101: oled_data = 16'b1111111111111111;
				14'b01101010110101: oled_data = 16'b1111111111111111;
				14'b01101100110101: oled_data = 16'b1111111111111111;
				14'b01101110110101: oled_data = 16'b1111111111111111;
				14'b01110000110101: oled_data = 16'b1111111111111111;
				14'b01110010110101: oled_data = 16'b1111111111111111;
				14'b01110100110101: oled_data = 16'b1111111111111111;
				14'b01110110110101: oled_data = 16'b1111111111111111;
				14'b01111000110101: oled_data = 16'b1111111111111111;
				14'b01111010110101: oled_data = 16'b1111111111111111;
				14'b01111100110101: oled_data = 16'b1111111111111111;
				14'b01111110110101: oled_data = 16'b1111111111111111;
				14'b10000000110101: oled_data = 16'b1111111111111111;
				14'b10000010110101: oled_data = 16'b1111111111111111;
				14'b10000100110101: oled_data = 16'b1111111111111111;
				14'b10000110110101: oled_data = 16'b1111111111111111;
				14'b10001000110101: oled_data = 16'b1111111111111111;
				14'b10001010110101: oled_data = 16'b1111111111111111;
				14'b10001100110101: oled_data = 16'b1111111111111111;
				14'b10001110110101: oled_data = 16'b1111111111111111;
				14'b10010000110101: oled_data = 16'b1111111111111111;
				14'b10010010110101: oled_data = 16'b1111111111111111;
				14'b10010100110101: oled_data = 16'b1111111111111111;
				14'b10010110110101: oled_data = 16'b1111111111111111;
				14'b10011000110101: oled_data = 16'b1111111111111111;
				14'b10011010110101: oled_data = 16'b1111111111111111;
				14'b10011100110101: oled_data = 16'b1111111111111111;
				14'b10011110110101: oled_data = 16'b1111111111111111;
				14'b10100000110101: oled_data = 16'b1111111111111111;
				14'b10100010110101: oled_data = 16'b1111111111111111;
				14'b10100100110101: oled_data = 16'b1111111111111111;
				14'b10100110110101: oled_data = 16'b1111111111111111;
				14'b10101000110101: oled_data = 16'b1111111111111111;
				14'b10101010110101: oled_data = 16'b1111111111111111;
				14'b10101100110101: oled_data = 16'b1111111111111111;
				14'b10101110110101: oled_data = 16'b1111111111111111;
				14'b10110000110101: oled_data = 16'b1111111111111111;
				14'b10110010110101: oled_data = 16'b1111111111111111;
				14'b10110100110101: oled_data = 16'b1111111111111111;
				14'b10110110110101: oled_data = 16'b1111111111111111;
				14'b10111000110101: oled_data = 16'b1111111111111111;
				14'b10111010110101: oled_data = 16'b1111111111111111;
				14'b10111100110101: oled_data = 16'b1111111111111111;
				14'b10111110110101: oled_data = 16'b1111111111111111;
				14'b00000000110110: oled_data = 16'b1111111111111111;
				14'b00000010110110: oled_data = 16'b1111111111111111;
				14'b00000100110110: oled_data = 16'b1111111111111111;
				14'b00000110110110: oled_data = 16'b1111111111111111;
				14'b00001000110110: oled_data = 16'b1111111111111111;
				14'b00001010110110: oled_data = 16'b1111111111111111;
				14'b00001100110110: oled_data = 16'b1111111111111111;
				14'b00001110110110: oled_data = 16'b1111111111111111;
				14'b00010000110110: oled_data = 16'b1111111111111111;
				14'b00010010110110: oled_data = 16'b1111111111111111;
				14'b00010100110110: oled_data = 16'b1111011110111110;
				14'b00010110110110: oled_data = 16'b1110011101111100;
				14'b00011000110110: oled_data = 16'b1101111101011011;
				14'b00011010110110: oled_data = 16'b1101011101011010;
				14'b00011100110110: oled_data = 16'b1100111100011001;
				14'b00011110110110: oled_data = 16'b1101111101111011;
				14'b00100000110110: oled_data = 16'b1111111111111110;
				14'b00100010110110: oled_data = 16'b1111111111111111;
				14'b00100100110110: oled_data = 16'b1111111111111111;
				14'b00100110110110: oled_data = 16'b1111111111111111;
				14'b00101000110110: oled_data = 16'b1111111111111111;
				14'b00101010110110: oled_data = 16'b1111111111111111;
				14'b00101100110110: oled_data = 16'b1111111111111111;
				14'b00101110110110: oled_data = 16'b1111111111111111;
				14'b00110000110110: oled_data = 16'b1111111111111111;
				14'b00110010110110: oled_data = 16'b1111111111111111;
				14'b00110100110110: oled_data = 16'b1111111111111111;
				14'b00110110110110: oled_data = 16'b1111111111111111;
				14'b00111000110110: oled_data = 16'b1111111111111111;
				14'b00111010110110: oled_data = 16'b1111111111111111;
				14'b00111100110110: oled_data = 16'b1111111111111111;
				14'b00111110110110: oled_data = 16'b1111111111111111;
				14'b01000000110110: oled_data = 16'b1111111111111111;
				14'b01000010110110: oled_data = 16'b1111111111111111;
				14'b01000100110110: oled_data = 16'b1111111111111111;
				14'b01000110110110: oled_data = 16'b1111111111111111;
				14'b01001000110110: oled_data = 16'b1111111111111111;
				14'b01001010110110: oled_data = 16'b1111111111111111;
				14'b01001100110110: oled_data = 16'b1111111111111111;
				14'b01001110110110: oled_data = 16'b1111111111111111;
				14'b01010000110110: oled_data = 16'b1111111111111111;
				14'b01010010110110: oled_data = 16'b1111111111111111;
				14'b01010100110110: oled_data = 16'b1111111111111111;
				14'b01010110110110: oled_data = 16'b1111111111111111;
				14'b01011000110110: oled_data = 16'b1111111111111111;
				14'b01011010110110: oled_data = 16'b1111111111111111;
				14'b01011100110110: oled_data = 16'b1111111111111111;
				14'b01011110110110: oled_data = 16'b1111111111111111;
				14'b01100000110110: oled_data = 16'b1111111111111111;
				14'b01100010110110: oled_data = 16'b1111111111111111;
				14'b01100100110110: oled_data = 16'b1111111111111111;
				14'b01100110110110: oled_data = 16'b1111111111111111;
				14'b01101000110110: oled_data = 16'b1111111111111111;
				14'b01101010110110: oled_data = 16'b1111111111111111;
				14'b01101100110110: oled_data = 16'b1111111111111111;
				14'b01101110110110: oled_data = 16'b1111111111111111;
				14'b01110000110110: oled_data = 16'b1111111111111111;
				14'b01110010110110: oled_data = 16'b1111111111111111;
				14'b01110100110110: oled_data = 16'b1111111111111111;
				14'b01110110110110: oled_data = 16'b1111111111111111;
				14'b01111000110110: oled_data = 16'b1111111111111111;
				14'b01111010110110: oled_data = 16'b1111111111111111;
				14'b01111100110110: oled_data = 16'b1111111111111111;
				14'b01111110110110: oled_data = 16'b1111111111111111;
				14'b10000000110110: oled_data = 16'b1111111111111111;
				14'b10000010110110: oled_data = 16'b1111111111111111;
				14'b10000100110110: oled_data = 16'b1111111111111111;
				14'b10000110110110: oled_data = 16'b1111111111111111;
				14'b10001000110110: oled_data = 16'b1111111111111111;
				14'b10001010110110: oled_data = 16'b1111111111111111;
				14'b10001100110110: oled_data = 16'b1111111111111111;
				14'b10001110110110: oled_data = 16'b1111111111111111;
				14'b10010000110110: oled_data = 16'b1111111111111111;
				14'b10010010110110: oled_data = 16'b1111111111111111;
				14'b10010100110110: oled_data = 16'b1111111111111111;
				14'b10010110110110: oled_data = 16'b1111111111111111;
				14'b10011000110110: oled_data = 16'b1111111111111111;
				14'b10011010110110: oled_data = 16'b1111111111111111;
				14'b10011100110110: oled_data = 16'b1111111111111111;
				14'b10011110110110: oled_data = 16'b1111111111111111;
				14'b10100000110110: oled_data = 16'b1111111111111111;
				14'b10100010110110: oled_data = 16'b1111111111111111;
				14'b10100100110110: oled_data = 16'b1111111111111111;
				14'b10100110110110: oled_data = 16'b1111111111111111;
				14'b10101000110110: oled_data = 16'b1111111111111111;
				14'b10101010110110: oled_data = 16'b1111111111111111;
				14'b10101100110110: oled_data = 16'b1111111111111111;
				14'b10101110110110: oled_data = 16'b1111111111111111;
				14'b10110000110110: oled_data = 16'b1111111111111111;
				14'b10110010110110: oled_data = 16'b1111111111111111;
				14'b10110100110110: oled_data = 16'b1111111111111111;
				14'b10110110110110: oled_data = 16'b1111111111111111;
				14'b10111000110110: oled_data = 16'b1111111111111111;
				14'b10111010110110: oled_data = 16'b1111111111111111;
				14'b10111100110110: oled_data = 16'b1111111111111111;
				14'b10111110110110: oled_data = 16'b1111111111111111;
				14'b00000000110111: oled_data = 16'b1111111111111111;
				14'b00000010110111: oled_data = 16'b1111111111111111;
				14'b00000100110111: oled_data = 16'b1111111111111111;
				14'b00000110110111: oled_data = 16'b1111111111111111;
				14'b00001000110111: oled_data = 16'b1111111111111111;
				14'b00001010110111: oled_data = 16'b1111111111111111;
				14'b00001100110111: oled_data = 16'b1111111111111111;
				14'b00001110110111: oled_data = 16'b1111111111111111;
				14'b00010000110111: oled_data = 16'b1111111111111111;
				14'b00010010110111: oled_data = 16'b1111111111111111;
				14'b00010100110111: oled_data = 16'b1111111111111111;
				14'b00010110110111: oled_data = 16'b1111011111011110;
				14'b00011000110111: oled_data = 16'b1110011101111100;
				14'b00011010110111: oled_data = 16'b1101111101011011;
				14'b00011100110111: oled_data = 16'b1101011101011010;
				14'b00011110110111: oled_data = 16'b1100111100011001;
				14'b00100000110111: oled_data = 16'b1110111110011100;
				14'b00100010110111: oled_data = 16'b1111111111111111;
				14'b00100100110111: oled_data = 16'b1111111111111111;
				14'b00100110110111: oled_data = 16'b1111111111111111;
				14'b00101000110111: oled_data = 16'b1111111111111111;
				14'b00101010110111: oled_data = 16'b1111111111111111;
				14'b00101100110111: oled_data = 16'b1111111111111111;
				14'b00101110110111: oled_data = 16'b1111111111111111;
				14'b00110000110111: oled_data = 16'b1111111111111111;
				14'b00110010110111: oled_data = 16'b1111111111111111;
				14'b00110100110111: oled_data = 16'b1111111111111111;
				14'b00110110110111: oled_data = 16'b1111111111111111;
				14'b00111000110111: oled_data = 16'b1111111111111111;
				14'b00111010110111: oled_data = 16'b1111111111111111;
				14'b00111100110111: oled_data = 16'b1111111111111111;
				14'b00111110110111: oled_data = 16'b1111111111111111;
				14'b01000000110111: oled_data = 16'b1111111111111111;
				14'b01000010110111: oled_data = 16'b1111111111111111;
				14'b01000100110111: oled_data = 16'b1111111111111111;
				14'b01000110110111: oled_data = 16'b1111111111111111;
				14'b01001000110111: oled_data = 16'b1111111111111111;
				14'b01001010110111: oled_data = 16'b1111111111111111;
				14'b01001100110111: oled_data = 16'b1111111111111111;
				14'b01001110110111: oled_data = 16'b1111111111111111;
				14'b01010000110111: oled_data = 16'b1111111111111111;
				14'b01010010110111: oled_data = 16'b1111111111111111;
				14'b01010100110111: oled_data = 16'b1111111111111111;
				14'b01010110110111: oled_data = 16'b1111111111111111;
				14'b01011000110111: oled_data = 16'b1111111111111111;
				14'b01011010110111: oled_data = 16'b1111111111111111;
				14'b01011100110111: oled_data = 16'b1111111111111111;
				14'b01011110110111: oled_data = 16'b1111111111111111;
				14'b01100000110111: oled_data = 16'b1111111111111111;
				14'b01100010110111: oled_data = 16'b1111111111111111;
				14'b01100100110111: oled_data = 16'b1111111111111111;
				14'b01100110110111: oled_data = 16'b1111111111111111;
				14'b01101000110111: oled_data = 16'b1111111111111111;
				14'b01101010110111: oled_data = 16'b1111111111111111;
				14'b01101100110111: oled_data = 16'b1111111111111111;
				14'b01101110110111: oled_data = 16'b1111111111111111;
				14'b01110000110111: oled_data = 16'b1111111111111111;
				14'b01110010110111: oled_data = 16'b1111111111111111;
				14'b01110100110111: oled_data = 16'b1111111111111111;
				14'b01110110110111: oled_data = 16'b1111111111111111;
				14'b01111000110111: oled_data = 16'b1111111111111111;
				14'b01111010110111: oled_data = 16'b1111111111111111;
				14'b01111100110111: oled_data = 16'b1111111111111111;
				14'b01111110110111: oled_data = 16'b1111111111111111;
				14'b10000000110111: oled_data = 16'b1111111111111111;
				14'b10000010110111: oled_data = 16'b1111111111111111;
				14'b10000100110111: oled_data = 16'b1111111111111111;
				14'b10000110110111: oled_data = 16'b1111111111111111;
				14'b10001000110111: oled_data = 16'b1111111111111111;
				14'b10001010110111: oled_data = 16'b1111111111111111;
				14'b10001100110111: oled_data = 16'b1111111111111111;
				14'b10001110110111: oled_data = 16'b1111111111111111;
				14'b10010000110111: oled_data = 16'b1111111111111111;
				14'b10010010110111: oled_data = 16'b1111111111111111;
				14'b10010100110111: oled_data = 16'b1111111111111111;
				14'b10010110110111: oled_data = 16'b1111111111111111;
				14'b10011000110111: oled_data = 16'b1111111111111111;
				14'b10011010110111: oled_data = 16'b1111111111111111;
				14'b10011100110111: oled_data = 16'b1111111111111111;
				14'b10011110110111: oled_data = 16'b1111111111111111;
				14'b10100000110111: oled_data = 16'b1111111111111111;
				14'b10100010110111: oled_data = 16'b1111111111111111;
				14'b10100100110111: oled_data = 16'b1111111111111111;
				14'b10100110110111: oled_data = 16'b1111111111111111;
				14'b10101000110111: oled_data = 16'b1111111111111111;
				14'b10101010110111: oled_data = 16'b1111111111111111;
				14'b10101100110111: oled_data = 16'b1111111111111111;
				14'b10101110110111: oled_data = 16'b1111111111111111;
				14'b10110000110111: oled_data = 16'b1111111111111111;
				14'b10110010110111: oled_data = 16'b1111111111111111;
				14'b10110100110111: oled_data = 16'b1111111111111111;
				14'b10110110110111: oled_data = 16'b1111111111111111;
				14'b10111000110111: oled_data = 16'b1111111111111111;
				14'b10111010110111: oled_data = 16'b1111111111111111;
				14'b10111100110111: oled_data = 16'b1111111111111111;
				14'b10111110110111: oled_data = 16'b1111111111111111;
				14'b00000000111000: oled_data = 16'b1111111111111111;
				14'b00000010111000: oled_data = 16'b1111111111111111;
				14'b00000100111000: oled_data = 16'b1111111111111111;
				14'b00000110111000: oled_data = 16'b1111111111111111;
				14'b00001000111000: oled_data = 16'b1111111111111111;
				14'b00001010111000: oled_data = 16'b1111111111111111;
				14'b00001100111000: oled_data = 16'b1111111111111111;
				14'b00001110111000: oled_data = 16'b1111111111111111;
				14'b00010000111000: oled_data = 16'b1111111111111111;
				14'b00010010111000: oled_data = 16'b1111111111111111;
				14'b00010100111000: oled_data = 16'b1111111111111111;
				14'b00010110111000: oled_data = 16'b1111111111111111;
				14'b00011000111000: oled_data = 16'b1111011111011110;
				14'b00011010111000: oled_data = 16'b1110011101111100;
				14'b00011100111000: oled_data = 16'b1101111101011011;
				14'b00011110111000: oled_data = 16'b1101011100111010;
				14'b00100000111000: oled_data = 16'b1101011100111001;
				14'b00100010111000: oled_data = 16'b1111011111011110;
				14'b00100100111000: oled_data = 16'b1111111111111111;
				14'b00100110111000: oled_data = 16'b1111111111111111;
				14'b00101000111000: oled_data = 16'b1111111111111111;
				14'b00101010111000: oled_data = 16'b1111111111111111;
				14'b00101100111000: oled_data = 16'b1111111111111111;
				14'b00101110111000: oled_data = 16'b1111111111111111;
				14'b00110000111000: oled_data = 16'b1111111111111111;
				14'b00110010111000: oled_data = 16'b1111111111111111;
				14'b00110100111000: oled_data = 16'b1111111111111111;
				14'b00110110111000: oled_data = 16'b1111111111111111;
				14'b00111000111000: oled_data = 16'b1111111111111111;
				14'b00111010111000: oled_data = 16'b1111111111111111;
				14'b00111100111000: oled_data = 16'b1111111111111111;
				14'b00111110111000: oled_data = 16'b1111111111111111;
				14'b01000000111000: oled_data = 16'b1111111111111111;
				14'b01000010111000: oled_data = 16'b1111111111111111;
				14'b01000100111000: oled_data = 16'b1111111111111111;
				14'b01000110111000: oled_data = 16'b1111111111111111;
				14'b01001000111000: oled_data = 16'b1111111111111111;
				14'b01001010111000: oled_data = 16'b1111111111111111;
				14'b01001100111000: oled_data = 16'b1111111111111111;
				14'b01001110111000: oled_data = 16'b1111111111111111;
				14'b01010000111000: oled_data = 16'b1111111111111111;
				14'b01010010111000: oled_data = 16'b1111111111111111;
				14'b01010100111000: oled_data = 16'b1111111111111111;
				14'b01010110111000: oled_data = 16'b1111111111111111;
				14'b01011000111000: oled_data = 16'b1111111111111111;
				14'b01011010111000: oled_data = 16'b1111111111111111;
				14'b01011100111000: oled_data = 16'b1111111111111111;
				14'b01011110111000: oled_data = 16'b1111111111111111;
				14'b01100000111000: oled_data = 16'b1111111111111111;
				14'b01100010111000: oled_data = 16'b1111111111111111;
				14'b01100100111000: oled_data = 16'b1111111111111111;
				14'b01100110111000: oled_data = 16'b1111111111111111;
				14'b01101000111000: oled_data = 16'b1111111111111111;
				14'b01101010111000: oled_data = 16'b1111111111111111;
				14'b01101100111000: oled_data = 16'b1111111111111111;
				14'b01101110111000: oled_data = 16'b1111111111111111;
				14'b01110000111000: oled_data = 16'b1111111111111111;
				14'b01110010111000: oled_data = 16'b1111111111111111;
				14'b01110100111000: oled_data = 16'b1111111111111111;
				14'b01110110111000: oled_data = 16'b1111111111111111;
				14'b01111000111000: oled_data = 16'b1111111111111111;
				14'b01111010111000: oled_data = 16'b1111111111111111;
				14'b01111100111000: oled_data = 16'b1111111111111111;
				14'b01111110111000: oled_data = 16'b1111111111111111;
				14'b10000000111000: oled_data = 16'b1111111111111111;
				14'b10000010111000: oled_data = 16'b1111111111111111;
				14'b10000100111000: oled_data = 16'b1111111111111111;
				14'b10000110111000: oled_data = 16'b1111111111111111;
				14'b10001000111000: oled_data = 16'b1111111111111111;
				14'b10001010111000: oled_data = 16'b1111111111111111;
				14'b10001100111000: oled_data = 16'b1111111111111111;
				14'b10001110111000: oled_data = 16'b1111111111111111;
				14'b10010000111000: oled_data = 16'b1111111111111111;
				14'b10010010111000: oled_data = 16'b1111111111111111;
				14'b10010100111000: oled_data = 16'b1111111111111111;
				14'b10010110111000: oled_data = 16'b1111111111111111;
				14'b10011000111000: oled_data = 16'b1111111111111111;
				14'b10011010111000: oled_data = 16'b1111111111111111;
				14'b10011100111000: oled_data = 16'b1111111111111111;
				14'b10011110111000: oled_data = 16'b1111111111111111;
				14'b10100000111000: oled_data = 16'b1111111111111111;
				14'b10100010111000: oled_data = 16'b1111111111111111;
				14'b10100100111000: oled_data = 16'b1111111111111111;
				14'b10100110111000: oled_data = 16'b1111111111111111;
				14'b10101000111000: oled_data = 16'b1111111111111111;
				14'b10101010111000: oled_data = 16'b1111111111111111;
				14'b10101100111000: oled_data = 16'b1111111111111111;
				14'b10101110111000: oled_data = 16'b1111111111111111;
				14'b10110000111000: oled_data = 16'b1111111111111111;
				14'b10110010111000: oled_data = 16'b1111111111111111;
				14'b10110100111000: oled_data = 16'b1111111111111111;
				14'b10110110111000: oled_data = 16'b1111111111111111;
				14'b10111000111000: oled_data = 16'b1111111111111111;
				14'b10111010111000: oled_data = 16'b1111111111111111;
				14'b10111100111000: oled_data = 16'b1111111111111111;
				14'b10111110111000: oled_data = 16'b1111111111111111;
				14'b00000000111001: oled_data = 16'b1111111111111111;
				14'b00000010111001: oled_data = 16'b1111111111111111;
				14'b00000100111001: oled_data = 16'b1111111111111111;
				14'b00000110111001: oled_data = 16'b1111111111111111;
				14'b00001000111001: oled_data = 16'b1111111111111111;
				14'b00001010111001: oled_data = 16'b1111111111111111;
				14'b00001100111001: oled_data = 16'b1111111111111111;
				14'b00001110111001: oled_data = 16'b1111111111111111;
				14'b00010000111001: oled_data = 16'b1111111111111111;
				14'b00010010111001: oled_data = 16'b1111111111111111;
				14'b00010100111001: oled_data = 16'b1111111111111111;
				14'b00010110111001: oled_data = 16'b1111111111111111;
				14'b00011000111001: oled_data = 16'b1111111111111111;
				14'b00011010111001: oled_data = 16'b1111011110111110;
				14'b00011100111001: oled_data = 16'b1101111101111011;
				14'b00011110111001: oled_data = 16'b1101111101011011;
				14'b00100000111001: oled_data = 16'b1101011100011001;
				14'b00100010111001: oled_data = 16'b1110011110011100;
				14'b00100100111001: oled_data = 16'b1111111111111111;
				14'b00100110111001: oled_data = 16'b1111111111111111;
				14'b00101000111001: oled_data = 16'b1111111111111111;
				14'b00101010111001: oled_data = 16'b1111111111111111;
				14'b00101100111001: oled_data = 16'b1111111111111111;
				14'b00101110111001: oled_data = 16'b1111111111111111;
				14'b00110000111001: oled_data = 16'b1111111111111111;
				14'b00110010111001: oled_data = 16'b1111111111111111;
				14'b00110100111001: oled_data = 16'b1111111111111111;
				14'b00110110111001: oled_data = 16'b1111111111111111;
				14'b00111000111001: oled_data = 16'b1111111111111111;
				14'b00111010111001: oled_data = 16'b1111111111111111;
				14'b00111100111001: oled_data = 16'b1111111111111111;
				14'b00111110111001: oled_data = 16'b1111111111111111;
				14'b01000000111001: oled_data = 16'b1111111111111111;
				14'b01000010111001: oled_data = 16'b1111111111111111;
				14'b01000100111001: oled_data = 16'b1111111111111111;
				14'b01000110111001: oled_data = 16'b1111111111111111;
				14'b01001000111001: oled_data = 16'b1111111111111111;
				14'b01001010111001: oled_data = 16'b1111111111111111;
				14'b01001100111001: oled_data = 16'b1111111111111111;
				14'b01001110111001: oled_data = 16'b1111111111111111;
				14'b01010000111001: oled_data = 16'b1111111111111111;
				14'b01010010111001: oled_data = 16'b1111111111111111;
				14'b01010100111001: oled_data = 16'b1111111111111111;
				14'b01010110111001: oled_data = 16'b1111111111111111;
				14'b01011000111001: oled_data = 16'b1111111111111111;
				14'b01011010111001: oled_data = 16'b1111111111111111;
				14'b01011100111001: oled_data = 16'b1111111111111111;
				14'b01011110111001: oled_data = 16'b1111111111111111;
				14'b01100000111001: oled_data = 16'b1111111111111111;
				14'b01100010111001: oled_data = 16'b1111111111111111;
				14'b01100100111001: oled_data = 16'b1111111111111111;
				14'b01100110111001: oled_data = 16'b1111111111111111;
				14'b01101000111001: oled_data = 16'b1111111111111111;
				14'b01101010111001: oled_data = 16'b1111111111111111;
				14'b01101100111001: oled_data = 16'b1111111111111111;
				14'b01101110111001: oled_data = 16'b1111111111111111;
				14'b01110000111001: oled_data = 16'b1111111111111111;
				14'b01110010111001: oled_data = 16'b1111111111111111;
				14'b01110100111001: oled_data = 16'b1111111111111111;
				14'b01110110111001: oled_data = 16'b1111111111111111;
				14'b01111000111001: oled_data = 16'b1111111111111111;
				14'b01111010111001: oled_data = 16'b1111111111111111;
				14'b01111100111001: oled_data = 16'b1111111111111111;
				14'b01111110111001: oled_data = 16'b1111111111111111;
				14'b10000000111001: oled_data = 16'b1111111111111111;
				14'b10000010111001: oled_data = 16'b1111111111111111;
				14'b10000100111001: oled_data = 16'b1111111111111111;
				14'b10000110111001: oled_data = 16'b1111111111111111;
				14'b10001000111001: oled_data = 16'b1111111111111111;
				14'b10001010111001: oled_data = 16'b1111111111111111;
				14'b10001100111001: oled_data = 16'b1111111111111111;
				14'b10001110111001: oled_data = 16'b1111111111111111;
				14'b10010000111001: oled_data = 16'b1111111111111111;
				14'b10010010111001: oled_data = 16'b1111111111111111;
				14'b10010100111001: oled_data = 16'b1111111111111111;
				14'b10010110111001: oled_data = 16'b1111111111111111;
				14'b10011000111001: oled_data = 16'b1111111111111111;
				14'b10011010111001: oled_data = 16'b1111111111111111;
				14'b10011100111001: oled_data = 16'b1111111111111111;
				14'b10011110111001: oled_data = 16'b1111111111111111;
				14'b10100000111001: oled_data = 16'b1111111111111111;
				14'b10100010111001: oled_data = 16'b1111111111111111;
				14'b10100100111001: oled_data = 16'b1111111111111111;
				14'b10100110111001: oled_data = 16'b1111111111111111;
				14'b10101000111001: oled_data = 16'b1111111111111111;
				14'b10101010111001: oled_data = 16'b1111111111111111;
				14'b10101100111001: oled_data = 16'b1111111111111111;
				14'b10101110111001: oled_data = 16'b1111111111111111;
				14'b10110000111001: oled_data = 16'b1111111111111111;
				14'b10110010111001: oled_data = 16'b1111111111111111;
				14'b10110100111001: oled_data = 16'b1111111111111111;
				14'b10110110111001: oled_data = 16'b1111111111111111;
				14'b10111000111001: oled_data = 16'b1111111111111111;
				14'b10111010111001: oled_data = 16'b1111111111111111;
				14'b10111100111001: oled_data = 16'b1111111111111111;
				14'b10111110111001: oled_data = 16'b1111111111111111;
				14'b00000000111010: oled_data = 16'b1111111111111111;
				14'b00000010111010: oled_data = 16'b1111111111111111;
				14'b00000100111010: oled_data = 16'b1111111111111111;
				14'b00000110111010: oled_data = 16'b1111111111111111;
				14'b00001000111010: oled_data = 16'b1111111111111111;
				14'b00001010111010: oled_data = 16'b1111111111111111;
				14'b00001100111010: oled_data = 16'b1111111111111111;
				14'b00001110111010: oled_data = 16'b1111111111111111;
				14'b00010000111010: oled_data = 16'b1111111111111111;
				14'b00010010111010: oled_data = 16'b1111111111111111;
				14'b00010100111010: oled_data = 16'b1111111111111111;
				14'b00010110111010: oled_data = 16'b1111111111111111;
				14'b00011000111010: oled_data = 16'b1111111111111111;
				14'b00011010111010: oled_data = 16'b1111111111111111;
				14'b00011100111010: oled_data = 16'b1110111110011101;
				14'b00011110111010: oled_data = 16'b1101111101011011;
				14'b00100000111010: oled_data = 16'b1101011100111010;
				14'b00100010111010: oled_data = 16'b1101011100111001;
				14'b00100100111010: oled_data = 16'b1111011111011110;
				14'b00100110111010: oled_data = 16'b1111111111111111;
				14'b00101000111010: oled_data = 16'b1111111111111111;
				14'b00101010111010: oled_data = 16'b1111111111111111;
				14'b00101100111010: oled_data = 16'b1111111111111111;
				14'b00101110111010: oled_data = 16'b1111111111111111;
				14'b00110000111010: oled_data = 16'b1111111111111111;
				14'b00110010111010: oled_data = 16'b1111111111111111;
				14'b00110100111010: oled_data = 16'b1111111111111111;
				14'b00110110111010: oled_data = 16'b1111111111111111;
				14'b00111000111010: oled_data = 16'b1111111111111111;
				14'b00111010111010: oled_data = 16'b1111111111111111;
				14'b00111100111010: oled_data = 16'b1111111111111111;
				14'b00111110111010: oled_data = 16'b1111111111111111;
				14'b01000000111010: oled_data = 16'b1111111111111111;
				14'b01000010111010: oled_data = 16'b1111111111111111;
				14'b01000100111010: oled_data = 16'b1111111111111111;
				14'b01000110111010: oled_data = 16'b1111111111111111;
				14'b01001000111010: oled_data = 16'b1111111111111111;
				14'b01001010111010: oled_data = 16'b1111111111111111;
				14'b01001100111010: oled_data = 16'b1111111111111111;
				14'b01001110111010: oled_data = 16'b1111111111111111;
				14'b01010000111010: oled_data = 16'b1111111111111111;
				14'b01010010111010: oled_data = 16'b1111111111111111;
				14'b01010100111010: oled_data = 16'b1111111111111111;
				14'b01010110111010: oled_data = 16'b1111111111111111;
				14'b01011000111010: oled_data = 16'b1111111111111111;
				14'b01011010111010: oled_data = 16'b1111111111111111;
				14'b01011100111010: oled_data = 16'b1111111111111111;
				14'b01011110111010: oled_data = 16'b1111111111111111;
				14'b01100000111010: oled_data = 16'b1111111111111111;
				14'b01100010111010: oled_data = 16'b1111111111111111;
				14'b01100100111010: oled_data = 16'b1111111111111111;
				14'b01100110111010: oled_data = 16'b1111111111111111;
				14'b01101000111010: oled_data = 16'b1111111111111111;
				14'b01101010111010: oled_data = 16'b1111111111111111;
				14'b01101100111010: oled_data = 16'b1111111111111111;
				14'b01101110111010: oled_data = 16'b1111111111111111;
				14'b01110000111010: oled_data = 16'b1111111111111111;
				14'b01110010111010: oled_data = 16'b1111111111111111;
				14'b01110100111010: oled_data = 16'b1111111111111111;
				14'b01110110111010: oled_data = 16'b1111111111111111;
				14'b01111000111010: oled_data = 16'b1111111111111111;
				14'b01111010111010: oled_data = 16'b1111111111111111;
				14'b01111100111010: oled_data = 16'b1111111111111111;
				14'b01111110111010: oled_data = 16'b1111111111111111;
				14'b10000000111010: oled_data = 16'b1111111111111111;
				14'b10000010111010: oled_data = 16'b1111111111111111;
				14'b10000100111010: oled_data = 16'b1111111111111111;
				14'b10000110111010: oled_data = 16'b1111111111111111;
				14'b10001000111010: oled_data = 16'b1111111111111111;
				14'b10001010111010: oled_data = 16'b1111111111111111;
				14'b10001100111010: oled_data = 16'b1111111111111111;
				14'b10001110111010: oled_data = 16'b1111111111111111;
				14'b10010000111010: oled_data = 16'b1111111111111111;
				14'b10010010111010: oled_data = 16'b1111111111111111;
				14'b10010100111010: oled_data = 16'b1111111111111111;
				14'b10010110111010: oled_data = 16'b1111111111111111;
				14'b10011000111010: oled_data = 16'b1111111111111111;
				14'b10011010111010: oled_data = 16'b1111111111111111;
				14'b10011100111010: oled_data = 16'b1111111111111111;
				14'b10011110111010: oled_data = 16'b1111111111111111;
				14'b10100000111010: oled_data = 16'b1111111111111111;
				14'b10100010111010: oled_data = 16'b1111111111111111;
				14'b10100100111010: oled_data = 16'b1111111111111111;
				14'b10100110111010: oled_data = 16'b1111111111111111;
				14'b10101000111010: oled_data = 16'b1111111111111111;
				14'b10101010111010: oled_data = 16'b1111111111111111;
				14'b10101100111010: oled_data = 16'b1111111111111111;
				14'b10101110111010: oled_data = 16'b1111111111111111;
				14'b10110000111010: oled_data = 16'b1111111111111111;
				14'b10110010111010: oled_data = 16'b1111111111111111;
				14'b10110100111010: oled_data = 16'b1111111111111111;
				14'b10110110111010: oled_data = 16'b1111111111111111;
				14'b10111000111010: oled_data = 16'b1111111111111111;
				14'b10111010111010: oled_data = 16'b1111111111111111;
				14'b10111100111010: oled_data = 16'b1111111111111111;
				14'b10111110111010: oled_data = 16'b1111111111111111;
				14'b00000000111011: oled_data = 16'b1111111111111111;
				14'b00000010111011: oled_data = 16'b1111111111111111;
				14'b00000100111011: oled_data = 16'b1111111111111111;
				14'b00000110111011: oled_data = 16'b1111111111111111;
				14'b00001000111011: oled_data = 16'b1111111111111111;
				14'b00001010111011: oled_data = 16'b1111111111111111;
				14'b00001100111011: oled_data = 16'b1111111111111111;
				14'b00001110111011: oled_data = 16'b1111111111111111;
				14'b00010000111011: oled_data = 16'b1111111111111111;
				14'b00010010111011: oled_data = 16'b1111111111111111;
				14'b00010100111011: oled_data = 16'b1111111111111111;
				14'b00010110111011: oled_data = 16'b1111111111111111;
				14'b00011000111011: oled_data = 16'b1111111111111111;
				14'b00011010111011: oled_data = 16'b1111111111111111;
				14'b00011100111011: oled_data = 16'b1111011111011110;
				14'b00011110111011: oled_data = 16'b1110011101111011;
				14'b00100000111011: oled_data = 16'b1101111101011010;
				14'b00100010111011: oled_data = 16'b1101011100111001;
				14'b00100100111011: oled_data = 16'b1110111110111101;
				14'b00100110111011: oled_data = 16'b1111111111111111;
				14'b00101000111011: oled_data = 16'b1111111111111111;
				14'b00101010111011: oled_data = 16'b1111111111111111;
				14'b00101100111011: oled_data = 16'b1111111111111111;
				14'b00101110111011: oled_data = 16'b1111111111111111;
				14'b00110000111011: oled_data = 16'b1111111111111111;
				14'b00110010111011: oled_data = 16'b1111111111111111;
				14'b00110100111011: oled_data = 16'b1111111111111111;
				14'b00110110111011: oled_data = 16'b1111111111111111;
				14'b00111000111011: oled_data = 16'b1111111111111111;
				14'b00111010111011: oled_data = 16'b1111111111111111;
				14'b00111100111011: oled_data = 16'b1111111111111111;
				14'b00111110111011: oled_data = 16'b1111111111111111;
				14'b01000000111011: oled_data = 16'b1111111111111111;
				14'b01000010111011: oled_data = 16'b1111111111111111;
				14'b01000100111011: oled_data = 16'b1111111111111111;
				14'b01000110111011: oled_data = 16'b1111111111111111;
				14'b01001000111011: oled_data = 16'b1111111111111111;
				14'b01001010111011: oled_data = 16'b1111111111111111;
				14'b01001100111011: oled_data = 16'b1111111111111111;
				14'b01001110111011: oled_data = 16'b1111111111111111;
				14'b01010000111011: oled_data = 16'b1111111111111111;
				14'b01010010111011: oled_data = 16'b1111111111111111;
				14'b01010100111011: oled_data = 16'b1111111111111111;
				14'b01010110111011: oled_data = 16'b1111111111111111;
				14'b01011000111011: oled_data = 16'b1111111111111111;
				14'b01011010111011: oled_data = 16'b1111111111111111;
				14'b01011100111011: oled_data = 16'b1111111111111111;
				14'b01011110111011: oled_data = 16'b1111111111111111;
				14'b01100000111011: oled_data = 16'b1111111111111111;
				14'b01100010111011: oled_data = 16'b1111111111111111;
				14'b01100100111011: oled_data = 16'b1111111111111111;
				14'b01100110111011: oled_data = 16'b1111111111111111;
				14'b01101000111011: oled_data = 16'b1111111111111111;
				14'b01101010111011: oled_data = 16'b1111111111111111;
				14'b01101100111011: oled_data = 16'b1111111111111111;
				14'b01101110111011: oled_data = 16'b1111111111111111;
				14'b01110000111011: oled_data = 16'b1111111111111111;
				14'b01110010111011: oled_data = 16'b1111111111111111;
				14'b01110100111011: oled_data = 16'b1111111111111111;
				14'b01110110111011: oled_data = 16'b1111111111111111;
				14'b01111000111011: oled_data = 16'b1111111111111111;
				14'b01111010111011: oled_data = 16'b1111111111111111;
				14'b01111100111011: oled_data = 16'b1111111111111111;
				14'b01111110111011: oled_data = 16'b1111111111111111;
				14'b10000000111011: oled_data = 16'b1111111111111111;
				14'b10000010111011: oled_data = 16'b1111111111111111;
				14'b10000100111011: oled_data = 16'b1111111111111111;
				14'b10000110111011: oled_data = 16'b1111111111111111;
				14'b10001000111011: oled_data = 16'b1111111111111111;
				14'b10001010111011: oled_data = 16'b1111111111111111;
				14'b10001100111011: oled_data = 16'b1111111111111111;
				14'b10001110111011: oled_data = 16'b1111111111111111;
				14'b10010000111011: oled_data = 16'b1111111111111111;
				14'b10010010111011: oled_data = 16'b1111111111111111;
				14'b10010100111011: oled_data = 16'b1111111111111111;
				14'b10010110111011: oled_data = 16'b1111111111111111;
				14'b10011000111011: oled_data = 16'b1111111111111111;
				14'b10011010111011: oled_data = 16'b1111111111111111;
				14'b10011100111011: oled_data = 16'b1111111111111111;
				14'b10011110111011: oled_data = 16'b1111111111111111;
				14'b10100000111011: oled_data = 16'b1111111111111111;
				14'b10100010111011: oled_data = 16'b1111111111111111;
				14'b10100100111011: oled_data = 16'b1111111111111111;
				14'b10100110111011: oled_data = 16'b1111111111111111;
				14'b10101000111011: oled_data = 16'b1111111111111111;
				14'b10101010111011: oled_data = 16'b1111111111111111;
				14'b10101100111011: oled_data = 16'b1111111111111111;
				14'b10101110111011: oled_data = 16'b1111111111111111;
				14'b10110000111011: oled_data = 16'b1111111111111111;
				14'b10110010111011: oled_data = 16'b1111111111111111;
				14'b10110100111011: oled_data = 16'b1111111111111111;
				14'b10110110111011: oled_data = 16'b1111111111111111;
				14'b10111000111011: oled_data = 16'b1111111111111111;
				14'b10111010111011: oled_data = 16'b1111111111111111;
				14'b10111100111011: oled_data = 16'b1111111111111111;
				14'b10111110111011: oled_data = 16'b1111111111111111;
				14'b00000000111100: oled_data = 16'b1111111111111111;
				14'b00000010111100: oled_data = 16'b1111111111111111;
				14'b00000100111100: oled_data = 16'b1111111111111111;
				14'b00000110111100: oled_data = 16'b1111111111111111;
				14'b00001000111100: oled_data = 16'b1111111111111111;
				14'b00001010111100: oled_data = 16'b1111111111111111;
				14'b00001100111100: oled_data = 16'b1111111111111111;
				14'b00001110111100: oled_data = 16'b1111111111111111;
				14'b00010000111100: oled_data = 16'b1111111111111111;
				14'b00010010111100: oled_data = 16'b1111111111111111;
				14'b00010100111100: oled_data = 16'b1111111111111111;
				14'b00010110111100: oled_data = 16'b1111111111111111;
				14'b00011000111100: oled_data = 16'b1111111111111111;
				14'b00011010111100: oled_data = 16'b1111111111111111;
				14'b00011100111100: oled_data = 16'b1111111111111111;
				14'b00011110111100: oled_data = 16'b1110111110011101;
				14'b00100000111100: oled_data = 16'b1101111101011011;
				14'b00100010111100: oled_data = 16'b1101011100111001;
				14'b00100100111100: oled_data = 16'b1110011101111011;
				14'b00100110111100: oled_data = 16'b1111111111111111;
				14'b00101000111100: oled_data = 16'b1111111111111111;
				14'b00101010111100: oled_data = 16'b1111111111111111;
				14'b00101100111100: oled_data = 16'b1111111111111111;
				14'b00101110111100: oled_data = 16'b1111111111111111;
				14'b00110000111100: oled_data = 16'b1111111111111111;
				14'b00110010111100: oled_data = 16'b1111111111111111;
				14'b00110100111100: oled_data = 16'b1111111111111111;
				14'b00110110111100: oled_data = 16'b1111111111111111;
				14'b00111000111100: oled_data = 16'b1111111111111111;
				14'b00111010111100: oled_data = 16'b1111111111111111;
				14'b00111100111100: oled_data = 16'b1111111111111111;
				14'b00111110111100: oled_data = 16'b1111111111111111;
				14'b01000000111100: oled_data = 16'b1111111111111111;
				14'b01000010111100: oled_data = 16'b1111111111111111;
				14'b01000100111100: oled_data = 16'b1111111111111111;
				14'b01000110111100: oled_data = 16'b1111111111111111;
				14'b01001000111100: oled_data = 16'b1111111111111111;
				14'b01001010111100: oled_data = 16'b1111111111111111;
				14'b01001100111100: oled_data = 16'b1111111111111111;
				14'b01001110111100: oled_data = 16'b1111111111111111;
				14'b01010000111100: oled_data = 16'b1111111111111111;
				14'b01010010111100: oled_data = 16'b1111111111111111;
				14'b01010100111100: oled_data = 16'b1111111111111111;
				14'b01010110111100: oled_data = 16'b1111111111111111;
				14'b01011000111100: oled_data = 16'b1111111111111111;
				14'b01011010111100: oled_data = 16'b1111111111111111;
				14'b01011100111100: oled_data = 16'b1111111111111111;
				14'b01011110111100: oled_data = 16'b1111111111111111;
				14'b01100000111100: oled_data = 16'b1111111111111111;
				14'b01100010111100: oled_data = 16'b1111111111111111;
				14'b01100100111100: oled_data = 16'b1111111111111111;
				14'b01100110111100: oled_data = 16'b1111111111111111;
				14'b01101000111100: oled_data = 16'b1111111111111111;
				14'b01101010111100: oled_data = 16'b1111111111111111;
				14'b01101100111100: oled_data = 16'b1111111111111111;
				14'b01101110111100: oled_data = 16'b1111111111111111;
				14'b01110000111100: oled_data = 16'b1111111111111111;
				14'b01110010111100: oled_data = 16'b1111111111111111;
				14'b01110100111100: oled_data = 16'b1111111111111111;
				14'b01110110111100: oled_data = 16'b1111111111111111;
				14'b01111000111100: oled_data = 16'b1111111111111111;
				14'b01111010111100: oled_data = 16'b1111111111111111;
				14'b01111100111100: oled_data = 16'b1111111111111111;
				14'b01111110111100: oled_data = 16'b1111111111111111;
				14'b10000000111100: oled_data = 16'b1111111111111111;
				14'b10000010111100: oled_data = 16'b1111111111111111;
				14'b10000100111100: oled_data = 16'b1111111111111111;
				14'b10000110111100: oled_data = 16'b1111111111111111;
				14'b10001000111100: oled_data = 16'b1111111111111111;
				14'b10001010111100: oled_data = 16'b1111111111111111;
				14'b10001100111100: oled_data = 16'b1111111111111111;
				14'b10001110111100: oled_data = 16'b1111111111111111;
				14'b10010000111100: oled_data = 16'b1111111111111111;
				14'b10010010111100: oled_data = 16'b1111111111111111;
				14'b10010100111100: oled_data = 16'b1111111111111111;
				14'b10010110111100: oled_data = 16'b1111111111111111;
				14'b10011000111100: oled_data = 16'b1111111111111111;
				14'b10011010111100: oled_data = 16'b1111111111111111;
				14'b10011100111100: oled_data = 16'b1111111111111111;
				14'b10011110111100: oled_data = 16'b1111111111111111;
				14'b10100000111100: oled_data = 16'b1111111111111111;
				14'b10100010111100: oled_data = 16'b1111111111111111;
				14'b10100100111100: oled_data = 16'b1111111111111111;
				14'b10100110111100: oled_data = 16'b1111111111111111;
				14'b10101000111100: oled_data = 16'b1111111111111111;
				14'b10101010111100: oled_data = 16'b1111111111111111;
				14'b10101100111100: oled_data = 16'b1111111111111111;
				14'b10101110111100: oled_data = 16'b1111111111111111;
				14'b10110000111100: oled_data = 16'b1111111111111111;
				14'b10110010111100: oled_data = 16'b1111111111111111;
				14'b10110100111100: oled_data = 16'b1111111111111111;
				14'b10110110111100: oled_data = 16'b1111111111111111;
				14'b10111000111100: oled_data = 16'b1111111111111111;
				14'b10111010111100: oled_data = 16'b1111111111111111;
				14'b10111100111100: oled_data = 16'b1111111111111111;
				14'b10111110111100: oled_data = 16'b1111111111111111;
				14'b00000000111101: oled_data = 16'b1111111111111111;
				14'b00000010111101: oled_data = 16'b1111111111111111;
				14'b00000100111101: oled_data = 16'b1111111111111111;
				14'b00000110111101: oled_data = 16'b1111111111111111;
				14'b00001000111101: oled_data = 16'b1111111111111111;
				14'b00001010111101: oled_data = 16'b1111111111111111;
				14'b00001100111101: oled_data = 16'b1111111111111111;
				14'b00001110111101: oled_data = 16'b1111111111111111;
				14'b00010000111101: oled_data = 16'b1111111111111111;
				14'b00010010111101: oled_data = 16'b1111111111111111;
				14'b00010100111101: oled_data = 16'b1111111111111111;
				14'b00010110111101: oled_data = 16'b1111111111111111;
				14'b00011000111101: oled_data = 16'b1111111111111111;
				14'b00011010111101: oled_data = 16'b1111111111111111;
				14'b00011100111101: oled_data = 16'b1111111111111111;
				14'b00011110111101: oled_data = 16'b1111011110111110;
				14'b00100000111101: oled_data = 16'b1101111101011011;
				14'b00100010111101: oled_data = 16'b1101011101011010;
				14'b00100100111101: oled_data = 16'b1101111101011010;
				14'b00100110111101: oled_data = 16'b1111111111111111;
				14'b00101000111101: oled_data = 16'b1111111111111111;
				14'b00101010111101: oled_data = 16'b1111111111111111;
				14'b00101100111101: oled_data = 16'b1111111111111111;
				14'b00101110111101: oled_data = 16'b1111111111111111;
				14'b00110000111101: oled_data = 16'b1111111111111111;
				14'b00110010111101: oled_data = 16'b1111111111111111;
				14'b00110100111101: oled_data = 16'b1111111111111111;
				14'b00110110111101: oled_data = 16'b1111111111111111;
				14'b00111000111101: oled_data = 16'b1111111111111111;
				14'b00111010111101: oled_data = 16'b1111111111111111;
				14'b00111100111101: oled_data = 16'b1111111111111111;
				14'b00111110111101: oled_data = 16'b1111111111111111;
				14'b01000000111101: oled_data = 16'b1111111111111111;
				14'b01000010111101: oled_data = 16'b1111111111111111;
				14'b01000100111101: oled_data = 16'b1111111111111111;
				14'b01000110111101: oled_data = 16'b1111111111111111;
				14'b01001000111101: oled_data = 16'b1111111111111111;
				14'b01001010111101: oled_data = 16'b1111111111111111;
				14'b01001100111101: oled_data = 16'b1111111111111111;
				14'b01001110111101: oled_data = 16'b1111111111111111;
				14'b01010000111101: oled_data = 16'b1111111111111111;
				14'b01010010111101: oled_data = 16'b1111111111111111;
				14'b01010100111101: oled_data = 16'b1111111111111111;
				14'b01010110111101: oled_data = 16'b1111111111111111;
				14'b01011000111101: oled_data = 16'b1111111111111111;
				14'b01011010111101: oled_data = 16'b1111111111111111;
				14'b01011100111101: oled_data = 16'b1111111111111111;
				14'b01011110111101: oled_data = 16'b1111111111111111;
				14'b01100000111101: oled_data = 16'b1111111111111111;
				14'b01100010111101: oled_data = 16'b1111111111111111;
				14'b01100100111101: oled_data = 16'b1111111111111111;
				14'b01100110111101: oled_data = 16'b1111111111111111;
				14'b01101000111101: oled_data = 16'b1111111111111111;
				14'b01101010111101: oled_data = 16'b1111111111111111;
				14'b01101100111101: oled_data = 16'b1111111111111111;
				14'b01101110111101: oled_data = 16'b1111111111111111;
				14'b01110000111101: oled_data = 16'b1111111111111111;
				14'b01110010111101: oled_data = 16'b1111111111111111;
				14'b01110100111101: oled_data = 16'b1111111111111111;
				14'b01110110111101: oled_data = 16'b1111111111111111;
				14'b01111000111101: oled_data = 16'b1111111111111111;
				14'b01111010111101: oled_data = 16'b1111111111111111;
				14'b01111100111101: oled_data = 16'b1111111111111111;
				14'b01111110111101: oled_data = 16'b1111111111111111;
				14'b10000000111101: oled_data = 16'b1111111111111111;
				14'b10000010111101: oled_data = 16'b1111111111111111;
				14'b10000100111101: oled_data = 16'b1111111111111111;
				14'b10000110111101: oled_data = 16'b1111111111111111;
				14'b10001000111101: oled_data = 16'b1111111111111111;
				14'b10001010111101: oled_data = 16'b1111111111111111;
				14'b10001100111101: oled_data = 16'b1111111111111111;
				14'b10001110111101: oled_data = 16'b1111111111111111;
				14'b10010000111101: oled_data = 16'b1111111111111111;
				14'b10010010111101: oled_data = 16'b1111111111111111;
				14'b10010100111101: oled_data = 16'b1111111111111111;
				14'b10010110111101: oled_data = 16'b1111111111111111;
				14'b10011000111101: oled_data = 16'b1111111111111111;
				14'b10011010111101: oled_data = 16'b1111111111111111;
				14'b10011100111101: oled_data = 16'b1111111111111111;
				14'b10011110111101: oled_data = 16'b1111111111111111;
				14'b10100000111101: oled_data = 16'b1111111111111111;
				14'b10100010111101: oled_data = 16'b1111111111111111;
				14'b10100100111101: oled_data = 16'b1111111111111111;
				14'b10100110111101: oled_data = 16'b1111111111111111;
				14'b10101000111101: oled_data = 16'b1111111111111111;
				14'b10101010111101: oled_data = 16'b1111111111111111;
				14'b10101100111101: oled_data = 16'b1111111111111111;
				14'b10101110111101: oled_data = 16'b1111111111111111;
				14'b10110000111101: oled_data = 16'b1111111111111111;
				14'b10110010111101: oled_data = 16'b1111111111111111;
				14'b10110100111101: oled_data = 16'b1111111111111111;
				14'b10110110111101: oled_data = 16'b1111111111111111;
				14'b10111000111101: oled_data = 16'b1111111111111111;
				14'b10111010111101: oled_data = 16'b1111111111111111;
				14'b10111100111101: oled_data = 16'b1111111111111111;
				14'b10111110111101: oled_data = 16'b1111111111111111;
				14'b00000000111110: oled_data = 16'b1111111111111111;
				14'b00000010111110: oled_data = 16'b1111111111111111;
				14'b00000100111110: oled_data = 16'b1111111111111111;
				14'b00000110111110: oled_data = 16'b1111111111111111;
				14'b00001000111110: oled_data = 16'b1111111111111111;
				14'b00001010111110: oled_data = 16'b1111111111111111;
				14'b00001100111110: oled_data = 16'b1111111111111111;
				14'b00001110111110: oled_data = 16'b1111111111111111;
				14'b00010000111110: oled_data = 16'b1111111111111111;
				14'b00010010111110: oled_data = 16'b1111111111111111;
				14'b00010100111110: oled_data = 16'b1111111111111111;
				14'b00010110111110: oled_data = 16'b1111111111111111;
				14'b00011000111110: oled_data = 16'b1111111111111111;
				14'b00011010111110: oled_data = 16'b1111111111111111;
				14'b00011100111110: oled_data = 16'b1111111111111111;
				14'b00011110111110: oled_data = 16'b1111011111011110;
				14'b00100000111110: oled_data = 16'b1101111101111011;
				14'b00100010111110: oled_data = 16'b1101111101011010;
				14'b00100100111110: oled_data = 16'b1101011101011010;
				14'b00100110111110: oled_data = 16'b1111011111011110;
				14'b00101000111110: oled_data = 16'b1111111111111111;
				14'b00101010111110: oled_data = 16'b1111111111111111;
				14'b00101100111110: oled_data = 16'b1111111111111111;
				14'b00101110111110: oled_data = 16'b1111111111111111;
				14'b00110000111110: oled_data = 16'b1111111111111111;
				14'b00110010111110: oled_data = 16'b1111111111111111;
				14'b00110100111110: oled_data = 16'b1111111111111111;
				14'b00110110111110: oled_data = 16'b1111111111111111;
				14'b00111000111110: oled_data = 16'b1111111111111111;
				14'b00111010111110: oled_data = 16'b1111111111111111;
				14'b00111100111110: oled_data = 16'b1111111111111111;
				14'b00111110111110: oled_data = 16'b1111111111111111;
				14'b01000000111110: oled_data = 16'b1111111111111111;
				14'b01000010111110: oled_data = 16'b1111111111111111;
				14'b01000100111110: oled_data = 16'b1111111111111111;
				14'b01000110111110: oled_data = 16'b1111111111111111;
				14'b01001000111110: oled_data = 16'b1111111111111111;
				14'b01001010111110: oled_data = 16'b1111111111111111;
				14'b01001100111110: oled_data = 16'b1111111111111111;
				14'b01001110111110: oled_data = 16'b1111111111111111;
				14'b01010000111110: oled_data = 16'b1111111111111111;
				14'b01010010111110: oled_data = 16'b1111111111111111;
				14'b01010100111110: oled_data = 16'b1111111111111111;
				14'b01010110111110: oled_data = 16'b1111111111111111;
				14'b01011000111110: oled_data = 16'b1111111111111111;
				14'b01011010111110: oled_data = 16'b1111111111111111;
				14'b01011100111110: oled_data = 16'b1111111111111111;
				14'b01011110111110: oled_data = 16'b1111111111111111;
				14'b01100000111110: oled_data = 16'b1111111111111111;
				14'b01100010111110: oled_data = 16'b1111111111111111;
				14'b01100100111110: oled_data = 16'b1111111111111111;
				14'b01100110111110: oled_data = 16'b1111111111111111;
				14'b01101000111110: oled_data = 16'b1111111111111111;
				14'b01101010111110: oled_data = 16'b1111111111111111;
				14'b01101100111110: oled_data = 16'b1111111111111111;
				14'b01101110111110: oled_data = 16'b1111111111111111;
				14'b01110000111110: oled_data = 16'b1111111111111111;
				14'b01110010111110: oled_data = 16'b1111111111111111;
				14'b01110100111110: oled_data = 16'b1111111111111111;
				14'b01110110111110: oled_data = 16'b1111111111111111;
				14'b01111000111110: oled_data = 16'b1111111111111111;
				14'b01111010111110: oled_data = 16'b1111111111111111;
				14'b01111100111110: oled_data = 16'b1111111111111111;
				14'b01111110111110: oled_data = 16'b1111111111111111;
				14'b10000000111110: oled_data = 16'b1111111111111111;
				14'b10000010111110: oled_data = 16'b1111111111111111;
				14'b10000100111110: oled_data = 16'b1111111111111111;
				14'b10000110111110: oled_data = 16'b1111111111111111;
				14'b10001000111110: oled_data = 16'b1111111111111111;
				14'b10001010111110: oled_data = 16'b1111111111111111;
				14'b10001100111110: oled_data = 16'b1111111111111111;
				14'b10001110111110: oled_data = 16'b1111111111111111;
				14'b10010000111110: oled_data = 16'b1111111111111111;
				14'b10010010111110: oled_data = 16'b1111111111111111;
				14'b10010100111110: oled_data = 16'b1111111111111111;
				14'b10010110111110: oled_data = 16'b1111111111111111;
				14'b10011000111110: oled_data = 16'b1111111111111111;
				14'b10011010111110: oled_data = 16'b1111111111111111;
				14'b10011100111110: oled_data = 16'b1111111111111111;
				14'b10011110111110: oled_data = 16'b1111111111111111;
				14'b10100000111110: oled_data = 16'b1111111111111111;
				14'b10100010111110: oled_data = 16'b1111111111111111;
				14'b10100100111110: oled_data = 16'b1111111111111111;
				14'b10100110111110: oled_data = 16'b1111111111111111;
				14'b10101000111110: oled_data = 16'b1111111111111111;
				14'b10101010111110: oled_data = 16'b1111111111111111;
				14'b10101100111110: oled_data = 16'b1111111111111111;
				14'b10101110111110: oled_data = 16'b1111111111111111;
				14'b10110000111110: oled_data = 16'b1111111111111111;
				14'b10110010111110: oled_data = 16'b1111111111111111;
				14'b10110100111110: oled_data = 16'b1111111111111111;
				14'b10110110111110: oled_data = 16'b1111111111111111;
				14'b10111000111110: oled_data = 16'b1111111111111111;
				14'b10111010111110: oled_data = 16'b1111111111111111;
				14'b10111100111110: oled_data = 16'b1111111111111111;
				14'b10111110111110: oled_data = 16'b1111111111111111;
				14'b00000000111111: oled_data = 16'b1111111111111111;
				14'b00000010111111: oled_data = 16'b1111111111111111;
				14'b00000100111111: oled_data = 16'b1111111111111111;
				14'b00000110111111: oled_data = 16'b1111111111111111;
				14'b00001000111111: oled_data = 16'b1111111111111111;
				14'b00001010111111: oled_data = 16'b1111111111111111;
				14'b00001100111111: oled_data = 16'b1111111111111111;
				14'b00001110111111: oled_data = 16'b1111111111111111;
				14'b00010000111111: oled_data = 16'b1111111111111111;
				14'b00010010111111: oled_data = 16'b1111111111111111;
				14'b00010100111111: oled_data = 16'b1111111111111111;
				14'b00010110111111: oled_data = 16'b1111111111111111;
				14'b00011000111111: oled_data = 16'b1111111111111111;
				14'b00011010111111: oled_data = 16'b1111111111111111;
				14'b00011100111111: oled_data = 16'b1111111111111111;
				14'b00011110111111: oled_data = 16'b1111011111011110;
				14'b00100000111111: oled_data = 16'b1110011101111100;
				14'b00100010111111: oled_data = 16'b1101111101011011;
				14'b00100100111111: oled_data = 16'b1101011100111010;
				14'b00100110111111: oled_data = 16'b1111011111011110;
				14'b00101000111111: oled_data = 16'b1111111111111111;
				14'b00101010111111: oled_data = 16'b1111111111111111;
				14'b00101100111111: oled_data = 16'b1111111111111111;
				14'b00101110111111: oled_data = 16'b1111111111111111;
				14'b00110000111111: oled_data = 16'b1111111111111111;
				14'b00110010111111: oled_data = 16'b1111111111111111;
				14'b00110100111111: oled_data = 16'b1111111111111111;
				14'b00110110111111: oled_data = 16'b1111111111111111;
				14'b00111000111111: oled_data = 16'b1111111111111111;
				14'b00111010111111: oled_data = 16'b1111111111111111;
				14'b00111100111111: oled_data = 16'b1111111111111111;
				14'b00111110111111: oled_data = 16'b1111111111111111;
				14'b01000000111111: oled_data = 16'b1111111111111111;
				14'b01000010111111: oled_data = 16'b1111111111111111;
				14'b01000100111111: oled_data = 16'b1111111111111111;
				14'b01000110111111: oled_data = 16'b1111111111111111;
				14'b01001000111111: oled_data = 16'b1111111111111111;
				14'b01001010111111: oled_data = 16'b1111111111111111;
				14'b01001100111111: oled_data = 16'b1111111111111111;
				14'b01001110111111: oled_data = 16'b1111111111111111;
				14'b01010000111111: oled_data = 16'b1111111111111111;
				14'b01010010111111: oled_data = 16'b1111111111111111;
				14'b01010100111111: oled_data = 16'b1111111111111111;
				14'b01010110111111: oled_data = 16'b1111111111111111;
				14'b01011000111111: oled_data = 16'b1111111111111111;
				14'b01011010111111: oled_data = 16'b1111111111111111;
				14'b01011100111111: oled_data = 16'b1111111111111111;
				14'b01011110111111: oled_data = 16'b1111111111111111;
				14'b01100000111111: oled_data = 16'b1111111111111111;
				14'b01100010111111: oled_data = 16'b1111111111111111;
				14'b01100100111111: oled_data = 16'b1111111111111111;
				14'b01100110111111: oled_data = 16'b1111111111111111;
				14'b01101000111111: oled_data = 16'b1111111111111111;
				14'b01101010111111: oled_data = 16'b1111111111111111;
				14'b01101100111111: oled_data = 16'b1111111111111111;
				14'b01101110111111: oled_data = 16'b1111111111111111;
				14'b01110000111111: oled_data = 16'b1111111111111111;
				14'b01110010111111: oled_data = 16'b1111111111111111;
				14'b01110100111111: oled_data = 16'b1111111111111111;
				14'b01110110111111: oled_data = 16'b1111111111111111;
				14'b01111000111111: oled_data = 16'b1111111111111111;
				14'b01111010111111: oled_data = 16'b1111111111111111;
				14'b01111100111111: oled_data = 16'b1111111111111111;
				14'b01111110111111: oled_data = 16'b1111111111111111;
				14'b10000000111111: oled_data = 16'b1111111111111111;
				14'b10000010111111: oled_data = 16'b1111111111111111;
				14'b10000100111111: oled_data = 16'b1111111111111111;
				14'b10000110111111: oled_data = 16'b1111111111111111;
				14'b10001000111111: oled_data = 16'b1111111111111111;
				14'b10001010111111: oled_data = 16'b1111111111111111;
				14'b10001100111111: oled_data = 16'b1111111111111111;
				14'b10001110111111: oled_data = 16'b1111111111111111;
				14'b10010000111111: oled_data = 16'b1111111111111111;
				14'b10010010111111: oled_data = 16'b1111111111111111;
				14'b10010100111111: oled_data = 16'b1111111111111111;
				14'b10010110111111: oled_data = 16'b1111111111111111;
				14'b10011000111111: oled_data = 16'b1111111111111111;
				14'b10011010111111: oled_data = 16'b1111111111111111;
				14'b10011100111111: oled_data = 16'b1111111111111111;
				14'b10011110111111: oled_data = 16'b1111111111111111;
				14'b10100000111111: oled_data = 16'b1111111111111111;
				14'b10100010111111: oled_data = 16'b1111111111111111;
				14'b10100100111111: oled_data = 16'b1111111111111111;
				14'b10100110111111: oled_data = 16'b1111111111111111;
				14'b10101000111111: oled_data = 16'b1111111111111111;
				14'b10101010111111: oled_data = 16'b1111111111111111;
				14'b10101100111111: oled_data = 16'b1111111111111111;
				14'b10101110111111: oled_data = 16'b1111111111111111;
				14'b10110000111111: oled_data = 16'b1111111111111111;
				14'b10110010111111: oled_data = 16'b1111111111111111;
				14'b10110100111111: oled_data = 16'b1111111111111111;
				14'b10110110111111: oled_data = 16'b1111111111111111;
				14'b10111000111111: oled_data = 16'b1111111111111111;
				14'b10111010111111: oled_data = 16'b1111111111111111;
				14'b10111100111111: oled_data = 16'b1111111111111111;
				14'b10111110111111: oled_data = 16'b1111111111111111;
			endcase

			case (menu_state)
				4'd1: if (sel1) oled_data = 16'b1111111111110101;
				4'd2: if (sel2) oled_data = 16'b1111111111110101;
				4'd3: if (sel3) oled_data = 16'b1111111111110101;
				4'd4: if (sel4) oled_data = 16'b1111111111110101;
				4'd5: if (sel5) oled_data = 16'b1111111111110101;
				4'd6: if (sel6) oled_data = 16'b1111111111110101;
				4'd7: if (sel7) oled_data = 16'b1111111111110101;
				4'd8: if (sel8) oled_data = 16'b1111111111110101;
				4'd9: if (sel9) oled_data = 16'b1111111111110101;
			endcase

			if (menu_state < 4'd6) begin
				case ({x, y})
					14'b00111110011010: oled_data = 16'b1111011100011001;
					14'b01000000011010: oled_data = 16'b1111011100011001;
					14'b01011100011010: oled_data = 16'b1110111101111101;
					14'b01011110011010: oled_data = 16'b1101111100011011;
					14'b01100000011010: oled_data = 16'b1101111100011011;
					14'b01100010011010: oled_data = 16'b1110111101111101;
					14'b00111100011011: oled_data = 16'b1111011010010110;
					14'b00111110011011: oled_data = 16'b1110001111000101;
					14'b01000000011011: oled_data = 16'b1110001111000110;
					14'b01000010011011: oled_data = 16'b1111011010110111;
					14'b01011000011011: oled_data = 16'b1110011101011100;
					14'b01011010011011: oled_data = 16'b1011110111110111;
					14'b01011100011011: oled_data = 16'b1011010110110110;
					14'b01011110011011: oled_data = 16'b1011110111110111;
					14'b01100000011011: oled_data = 16'b1011110111110111;
					14'b01100010011011: oled_data = 16'b1011010110110110;
					14'b01100100011011: oled_data = 16'b1011110111110111;
					14'b01100110011011: oled_data = 16'b1110011101011100;
					14'b00110100011100: oled_data = 16'b1111011101111100;
					14'b00110110011100: oled_data = 16'b1111011110111101;
					14'b00111100011100: oled_data = 16'b1110110110010000;
					14'b00111110011100: oled_data = 16'b1110001110000100;
					14'b01000000011100: oled_data = 16'b1110110011001100;
					14'b01000010011100: oled_data = 16'b1111011010010111;
					14'b01001000011100: oled_data = 16'b1111011110111101;
					14'b01001010011100: oled_data = 16'b1111011101111011;
					14'b01010110011100: oled_data = 16'b1101111100011011;
					14'b01011000011100: oled_data = 16'b1010110101110101;
					14'b01011010011100: oled_data = 16'b1101011011011010;
					14'b01011100011100: oled_data = 16'b1111011111011110;
					14'b01100010011100: oled_data = 16'b1111011111011110;
					14'b01100100011100: oled_data = 16'b1101011011011010;
					14'b01100110011100: oled_data = 16'b1010110101110101;
					14'b01101000011100: oled_data = 16'b1101111100011011;
					14'b01110110011100: oled_data = 16'b1111111101111000;
					14'b01111000011100: oled_data = 16'b1111111011001110;
					14'b01111010011100: oled_data = 16'b1111111100010010;
					14'b00110010011101: oled_data = 16'b1111111111011110;
					14'b00110100011101: oled_data = 16'b1110110110010000;
					14'b00110110011101: oled_data = 16'b1111011010010110;
					14'b00111000011101: oled_data = 16'b1111011110011101;
					14'b00111100011101: oled_data = 16'b1110110110110001;
					14'b00111110011101: oled_data = 16'b1110001110100100;
					14'b01000000011101: oled_data = 16'b1110110011001011;
					14'b01000010011101: oled_data = 16'b1111011010010110;
					14'b01000110011101: oled_data = 16'b1111011110011101;
					14'b01001000011101: oled_data = 16'b1111011010010110;
					14'b01001010011101: oled_data = 16'b1110110110010000;
					14'b01001100011101: oled_data = 16'b1111111111011110;
					14'b01010100011101: oled_data = 16'b1110111110011101;
					14'b01010110011101: oled_data = 16'b1010110101110101;
					14'b01011000011101: oled_data = 16'b1110011100111100;
					14'b01100110011101: oled_data = 16'b1110011100111100;
					14'b01101000011101: oled_data = 16'b1010110101110101;
					14'b01101010011101: oled_data = 16'b1110111110011101;
					14'b01110100011101: oled_data = 16'b1111111101010101;
					14'b01110110011101: oled_data = 16'b1111111011001100;
					14'b01111000011101: oled_data = 16'b1111111110011001;
					14'b01111010011101: oled_data = 16'b1111111111011110;
					14'b00110010011110: oled_data = 16'b1111011100011010;
					14'b00110100011110: oled_data = 16'b1110110110110001;
					14'b00110110011110: oled_data = 16'b1110110110010000;
					14'b00111000011110: oled_data = 16'b1111011110111101;
					14'b00111010011110: oled_data = 16'b1111111111011110;
					14'b00111100011110: oled_data = 16'b1110110110110001;
					14'b00111110011110: oled_data = 16'b1110001110100100;
					14'b01000000011110: oled_data = 16'b1110110011001011;
					14'b01000010011110: oled_data = 16'b1111011010010110;
					14'b01000100011110: oled_data = 16'b1111111111011110;
					14'b01000110011110: oled_data = 16'b1111011110111101;
					14'b01001000011110: oled_data = 16'b1110110110010000;
					14'b01001010011110: oled_data = 16'b1110110110110001;
					14'b01001100011110: oled_data = 16'b1111011100011010;
					14'b01010100011110: oled_data = 16'b1100111001011001;
					14'b01010110011110: oled_data = 16'b1100011001011000;
					14'b01101000011110: oled_data = 16'b1100011001011000;
					14'b01101010011110: oled_data = 16'b1100111001011001;
					14'b01110010011110: oled_data = 16'b1111111110111100;
					14'b01110100011110: oled_data = 16'b1111111010101011;
					14'b01110110011110: oled_data = 16'b1111111111011110;
					14'b01111010011110: oled_data = 16'b1111111110011000;
					14'b01111100011110: oled_data = 16'b1111111100010010;
					14'b01111110011110: oled_data = 16'b1111111100110100;
					14'b10000000011110: oled_data = 16'b1111111110111011;
					14'b10000010011110: oled_data = 16'b1111111111011100;
					14'b10000100011110: oled_data = 16'b1111111111011100;
					14'b00110010011111: oled_data = 16'b1111011011011000;
					14'b00110100011111: oled_data = 16'b1110110111010010;
					14'b00110110011111: oled_data = 16'b1111010111010010;
					14'b00111010011111: oled_data = 16'b1111010111010010;
					14'b00111100011111: oled_data = 16'b1110110101001110;
					14'b00111110011111: oled_data = 16'b1110001110100100;
					14'b01000000011111: oled_data = 16'b1110110011101100;
					14'b01000010011111: oled_data = 16'b1111011001010100;
					14'b01000100011111: oled_data = 16'b1111010111010010;
					14'b01001000011111: oled_data = 16'b1111010111010010;
					14'b01001010011111: oled_data = 16'b1110110111010010;
					14'b01001100011111: oled_data = 16'b1111011011011000;
					14'b01010010011111: oled_data = 16'b1111011111011110;
					14'b01010100011111: oled_data = 16'b1011010110110110;
					14'b01010110011111: oled_data = 16'b1110011101011100;
					14'b01101000011111: oled_data = 16'b1110011101011100;
					14'b01101010011111: oled_data = 16'b1011010110110110;
					14'b01101100011111: oled_data = 16'b1111011111011110;
					14'b01110010011111: oled_data = 16'b1111111101110111;
					14'b01110100011111: oled_data = 16'b1111111100010001;
					14'b01111000011111: oled_data = 16'b1111111011101111;
					14'b01111010011111: oled_data = 16'b1111110111100000;
					14'b01111100011111: oled_data = 16'b1111110111000000;
					14'b01111110011111: oled_data = 16'b1111110111000000;
					14'b10000000011111: oled_data = 16'b1111111000000010;
					14'b10000010011111: oled_data = 16'b1111111001100110;
					14'b10000100011111: oled_data = 16'b1111111001000101;
					14'b10000110011111: oled_data = 16'b1111111011101111;
					14'b10001000011111: oled_data = 16'b1111111101010100;
					14'b10001010011111: oled_data = 16'b1111111110011001;
					14'b10001100011111: oled_data = 16'b1111111111111110;
					14'b00110010100000: oled_data = 16'b1111011100111010;
					14'b00110100100000: oled_data = 16'b1110110110110001;
					14'b00110110100000: oled_data = 16'b1110110110110001;
					14'b00111000100000: oled_data = 16'b1111011110111101;
					14'b00111010100000: oled_data = 16'b1110110101101111;
					14'b00111100100000: oled_data = 16'b1110110101101111;
					14'b00111110100000: oled_data = 16'b1110001110000100;
					14'b01000000100000: oled_data = 16'b1110110001101001;
					14'b01000010100000: oled_data = 16'b1111011000010011;
					14'b01000100100000: oled_data = 16'b1110110101101111;
					14'b01000110100000: oled_data = 16'b1111011110111101;
					14'b01001000100000: oled_data = 16'b1110110110110001;
					14'b01001010100000: oled_data = 16'b1110110110110001;
					14'b01001100100000: oled_data = 16'b1111011100111010;
					14'b01010010100000: oled_data = 16'b1111011111011110;
					14'b01010100100000: oled_data = 16'b1011010110110110;
					14'b01010110100000: oled_data = 16'b1110011101011100;
					14'b01011000100000: oled_data = 16'b1101011011011010;
					14'b01011010100000: oled_data = 16'b1110011100111100;
					14'b01100100100000: oled_data = 16'b1110011100111100;
					14'b01100110100000: oled_data = 16'b1101011011011010;
					14'b01101000100000: oled_data = 16'b1110011101011100;
					14'b01101010100000: oled_data = 16'b1011010110110110;
					14'b01101100100000: oled_data = 16'b1111011111011110;
					14'b01110010100000: oled_data = 16'b1111111101110111;
					14'b01110100100000: oled_data = 16'b1111111100010010;
					14'b01110110100000: oled_data = 16'b1111111110011001;
					14'b01111000100000: oled_data = 16'b1111110111100000;
					14'b01111010100000: oled_data = 16'b1111110111100000;
					14'b01111100100000: oled_data = 16'b1111111000100011;
					14'b01111110100000: oled_data = 16'b1111110111100000;
					14'b10000000100000: oled_data = 16'b1111110111100000;
					14'b10000010100000: oled_data = 16'b1111110111100000;
					14'b10000100100000: oled_data = 16'b1111110111100000;
					14'b10000110100000: oled_data = 16'b1111110111000000;
					14'b10001000100000: oled_data = 16'b1111110111000000;
					14'b10001010100000: oled_data = 16'b1111111000100100;
					14'b10001100100000: oled_data = 16'b1111111110111100;
					14'b00110010100001: oled_data = 16'b1111111111011110;
					14'b00110100100001: oled_data = 16'b1110110110010000;
					14'b00110110100001: oled_data = 16'b1111011011011000;
					14'b00111000100001: oled_data = 16'b1111111111011110;
					14'b00111010100001: oled_data = 16'b1111011000010100;
					14'b00111100100001: oled_data = 16'b1110110101101111;
					14'b00111110100001: oled_data = 16'b1110110100001101;
					14'b01000000100001: oled_data = 16'b1110110100001101;
					14'b01000010100001: oled_data = 16'b1110110101001111;
					14'b01000100100001: oled_data = 16'b1111011000110100;
					14'b01000110100001: oled_data = 16'b1111011111011110;
					14'b01001000100001: oled_data = 16'b1111011011011000;
					14'b01001010100001: oled_data = 16'b1110110110010000;
					14'b01001100100001: oled_data = 16'b1111111111011110;
					14'b01010010100001: oled_data = 16'b1111011111011110;
					14'b01010100100001: oled_data = 16'b1011010111010110;
					14'b01010110100001: oled_data = 16'b1101011010111010;
					14'b01011000100001: oled_data = 16'b1001110011110011;
					14'b01011010100001: oled_data = 16'b1011010110010110;
					14'b01100100100001: oled_data = 16'b1011010110010110;
					14'b01100110100001: oled_data = 16'b1001110011110011;
					14'b01101000100001: oled_data = 16'b1101011010111010;
					14'b01101010100001: oled_data = 16'b1011010111010110;
					14'b01101100100001: oled_data = 16'b1111011111011110;
					14'b01110010100001: oled_data = 16'b1111111111011101;
					14'b01110100100001: oled_data = 16'b1111111011001101;
					14'b01110110100001: oled_data = 16'b1111111100010001;
					14'b01111000100001: oled_data = 16'b1111110111000000;
					14'b01111010100001: oled_data = 16'b1111110111100000;
					14'b01111100100001: oled_data = 16'b1111111011001101;
					14'b01111110100001: oled_data = 16'b1111111000100100;
					14'b10000000100001: oled_data = 16'b1111110111000000;
					14'b10000010100001: oled_data = 16'b1111110111100000;
					14'b10000100100001: oled_data = 16'b1111110111100000;
					14'b10000110100001: oled_data = 16'b1111110111100001;
					14'b10001000100001: oled_data = 16'b1111111010101100;
					14'b10001010100001: oled_data = 16'b1111111110011010;
					14'b00110100100010: oled_data = 16'b1111011110011100;
					14'b00110110100010: oled_data = 16'b1111011110111101;
					14'b00111010100010: oled_data = 16'b1111011110111110;
					14'b00111100100010: oled_data = 16'b1110110110110001;
					14'b00111110100010: oled_data = 16'b1110110100101110;
					14'b01000000100010: oled_data = 16'b1110110100101110;
					14'b01000010100010: oled_data = 16'b1110110111010001;
					14'b01000100100010: oled_data = 16'b1111011111011110;
					14'b01001000100010: oled_data = 16'b1111011110111101;
					14'b01001010100010: oled_data = 16'b1111011110011100;
					14'b01010010100010: oled_data = 16'b1111011111011110;
					14'b01010100100010: oled_data = 16'b1011010110010110;
					14'b01010110100010: oled_data = 16'b1011110111110111;
					14'b01011000100010: oled_data = 16'b1001110100010011;
					14'b01011010100010: oled_data = 16'b1011010110110110;
					14'b01100100100010: oled_data = 16'b1011010110110110;
					14'b01100110100010: oled_data = 16'b1001110100010011;
					14'b01101000100010: oled_data = 16'b1011110111110111;
					14'b01101010100010: oled_data = 16'b1011010110010110;
					14'b01101100100010: oled_data = 16'b1111011111011110;
					14'b01110100100010: oled_data = 16'b1111111101110111;
					14'b01110110100010: oled_data = 16'b1111111001100111;
					14'b01111000100010: oled_data = 16'b1111110111000000;
					14'b01111010100010: oled_data = 16'b1111110111000000;
					14'b01111100100010: oled_data = 16'b1111111001000110;
					14'b01111110100010: oled_data = 16'b1111111011101111;
					14'b10000000100010: oled_data = 16'b1111110111100000;
					14'b10000010100010: oled_data = 16'b1111110111000000;
					14'b10000100100010: oled_data = 16'b1111111000000001;
					14'b10000110100010: oled_data = 16'b1111111101010110;
					14'b00111110100011: oled_data = 16'b1111011000110100;
					14'b01000000100011: oled_data = 16'b1111011000110100;
					14'b01010010100011: oled_data = 16'b1111011111011110;
					14'b01010100100011: oled_data = 16'b1100011001011000;
					14'b01010110100011: oled_data = 16'b1100011001011000;
					14'b01011000100011: oled_data = 16'b1001110011110011;
					14'b01011010100011: oled_data = 16'b1011010110010110;
					14'b01100100100011: oled_data = 16'b1011010110110110;
					14'b01100110100011: oled_data = 16'b1001110011110011;
					14'b01101000100011: oled_data = 16'b1100011001011000;
					14'b01101010100011: oled_data = 16'b1100011001011000;
					14'b01101100100011: oled_data = 16'b1111011111011110;
					14'b01110110100011: oled_data = 16'b1111111110011010;
					14'b01111000100011: oled_data = 16'b1111111011101111;
					14'b01111010100011: oled_data = 16'b1111111010001010;
					14'b01111100100011: oled_data = 16'b1111111010001010;
					14'b01111110100011: oled_data = 16'b1111111100110011;
					14'b10000000100011: oled_data = 16'b1111111011110000;
					14'b10000010100011: oled_data = 16'b1111111010001010;
					14'b10000100100011: oled_data = 16'b1111111010001011;
					14'b10000110100011: oled_data = 16'b1111111110011010;
					14'b00111000100100: oled_data = 16'b1111111111011110;
					14'b00111010100100: oled_data = 16'b1111011000110100;
					14'b00111100100100: oled_data = 16'b1110110111010001;
					14'b00111110100100: oled_data = 16'b1110110100001101;
					14'b01000000100100: oled_data = 16'b1110110100001101;
					14'b01000010100100: oled_data = 16'b1110110111010001;
					14'b01000100100100: oled_data = 16'b1111011000110100;
					14'b01000110100100: oled_data = 16'b1111111111011110;
					14'b01010110100100: oled_data = 16'b1101111100011011;
					14'b01011000100100: oled_data = 16'b1001110011110011;
					14'b01011010100100: oled_data = 16'b1011010110110110;
					14'b01100100100100: oled_data = 16'b1011010110110110;
					14'b01100110100100: oled_data = 16'b1001110011110011;
					14'b01101000100100: oled_data = 16'b1101111100011011;
					14'b00111000100101: oled_data = 16'b1111111111111110;
					14'b00111010100101: oled_data = 16'b1111011100011001;
					14'b00111100100101: oled_data = 16'b1111011011011000;
					14'b00111110100101: oled_data = 16'b1111011011111001;
					14'b01000000100101: oled_data = 16'b1111011011111001;
					14'b01000010100101: oled_data = 16'b1111011011011000;
					14'b01000100100101: oled_data = 16'b1111011100011001;
					14'b01000110100101: oled_data = 16'b1111111111011110;
					14'b01010110100101: oled_data = 16'b1111011111011110;
					14'b01011000100101: oled_data = 16'b1110011100111100;
					14'b01011010100101: oled_data = 16'b1110111110011101;
					14'b01100100100101: oled_data = 16'b1110111110011101;
					14'b01100110100101: oled_data = 16'b1110011100111100;
					14'b01101000100101: oled_data = 16'b1111011111011110;
					14'b01000100101011: oled_data = 16'b1110011110011110;
					14'b01000110101011: oled_data = 16'b1101111101011110;
					14'b01001000101011: oled_data = 16'b1101111101011110;
					14'b01001010101011: oled_data = 16'b1101111101011110;
					14'b01001100101011: oled_data = 16'b1101111101011110;
					14'b01001110101011: oled_data = 16'b1101111101011110;
					14'b01010000101011: oled_data = 16'b1101111101011110;
					14'b01010010101011: oled_data = 16'b1101111101011110;
					14'b01010100101011: oled_data = 16'b1101111101011110;
					14'b01010110101011: oled_data = 16'b1101111101011110;
					14'b01011000101011: oled_data = 16'b1101111101011110;
					14'b01011010101011: oled_data = 16'b1101111101111110;
					14'b01011100101011: oled_data = 16'b1111011111011111;
					14'b01000010101100: oled_data = 16'b1110111110011110;
					14'b01000100101100: oled_data = 16'b0110110101011010;
					14'b01000110101100: oled_data = 16'b0111110110011011;
					14'b01001000101100: oled_data = 16'b1000010110011011;
					14'b01001010101100: oled_data = 16'b1000010110011011;
					14'b01001100101100: oled_data = 16'b1000010110011011;
					14'b01001110101100: oled_data = 16'b1000010110011011;
					14'b01010000101100: oled_data = 16'b1000010110011011;
					14'b01010010101100: oled_data = 16'b1000010110011011;
					14'b01010100101100: oled_data = 16'b1000010110011011;
					14'b01010110101100: oled_data = 16'b1000010110011011;
					14'b01011000101100: oled_data = 16'b1000010110011011;
					14'b01011010101100: oled_data = 16'b0110110100111010;
					14'b01011100101100: oled_data = 16'b1100111100011101;
					14'b01100100101100: oled_data = 16'b1111011111011110;
					14'b01100110101100: oled_data = 16'b1101111101011010;
					14'b01101000101100: oled_data = 16'b1101011100111001;
					14'b01101010101100: oled_data = 16'b1101011100111001;
					14'b01101100101100: oled_data = 16'b1101011100111001;
					14'b01101110101100: oled_data = 16'b1101011100111001;
					14'b01110000101100: oled_data = 16'b1101011100111001;
					14'b01110010101100: oled_data = 16'b1101011100111001;
					14'b01110100101100: oled_data = 16'b1101011100111001;
					14'b01110110101100: oled_data = 16'b1101011100111001;
					14'b01111000101100: oled_data = 16'b1101111101011010;
					14'b01111010101100: oled_data = 16'b1111011111011110;
					14'b01000010101101: oled_data = 16'b1110011101111110;
					14'b01000100101101: oled_data = 16'b0111110101111011;
					14'b01000110101101: oled_data = 16'b1111011111011110;
					14'b01011010101101: oled_data = 16'b1000110111011011;
					14'b01011100101101: oled_data = 16'b1100011011011101;
					14'b01100100101101: oled_data = 16'b1101011101011001;
					14'b01100110101101: oled_data = 16'b0111110110001010;
					14'b01101000101101: oled_data = 16'b1001011000001110;
					14'b01101010101101: oled_data = 16'b1001011000001110;
					14'b01101100101101: oled_data = 16'b1001011000001110;
					14'b01101110101101: oled_data = 16'b1001011000001110;
					14'b01110000101101: oled_data = 16'b1001011000001110;
					14'b01110010101101: oled_data = 16'b1001011000001110;
					14'b01110100101101: oled_data = 16'b1001011000001110;
					14'b01110110101101: oled_data = 16'b1001011000001110;
					14'b01111000101101: oled_data = 16'b0111110110001010;
					14'b01111010101101: oled_data = 16'b1101011101011001;
					14'b01000010101110: oled_data = 16'b1110011101111110;
					14'b01000100101110: oled_data = 16'b0111110101111011;
					14'b01000110101110: oled_data = 16'b1111011111011110;
					14'b01011010101110: oled_data = 16'b1000110111011011;
					14'b01011100101110: oled_data = 16'b1100011011011101;
					14'b01100100101110: oled_data = 16'b1100111100011000;
					14'b01100110101110: oled_data = 16'b1001111000101111;
					14'b01111000101110: oled_data = 16'b1001111000101111;
					14'b01111010101110: oled_data = 16'b1100111100111000;
					14'b01000010101111: oled_data = 16'b1110011101111110;
					14'b01000100101111: oled_data = 16'b0111110101111011;
					14'b01000110101111: oled_data = 16'b1111011111011110;
					14'b01011010101111: oled_data = 16'b1000110111011011;
					14'b01011100101111: oled_data = 16'b1100011011011101;
					14'b01100100101111: oled_data = 16'b1100111100011000;
					14'b01100110101111: oled_data = 16'b1001111000101111;
					14'b01111000101111: oled_data = 16'b1001111000101111;
					14'b01111010101111: oled_data = 16'b1100111100111000;
					14'b01000010110000: oled_data = 16'b1110011101111110;
					14'b01000100110000: oled_data = 16'b0111110101111011;
					14'b01000110110000: oled_data = 16'b1111011111011110;
					14'b01011010110000: oled_data = 16'b1000110111011011;
					14'b01011100110000: oled_data = 16'b1100011011011101;
					14'b01100100110000: oled_data = 16'b1100111100011000;
					14'b01100110110000: oled_data = 16'b1001111000101111;
					14'b01111000110000: oled_data = 16'b1001111000101111;
					14'b01111010110000: oled_data = 16'b1100111100111000;
					14'b01000010110001: oled_data = 16'b1110011101111110;
					14'b01000100110001: oled_data = 16'b0111110101111011;
					14'b01000110110001: oled_data = 16'b1111011111011110;
					14'b01011010110001: oled_data = 16'b1000110111011011;
					14'b01011100110001: oled_data = 16'b1100011011011101;
					14'b01100100110001: oled_data = 16'b1100111100011000;
					14'b01100110110001: oled_data = 16'b1001111000101111;
					14'b01111000110001: oled_data = 16'b1001111000101111;
					14'b01111010110001: oled_data = 16'b1100111100111000;
					14'b01000010110010: oled_data = 16'b1110011101111110;
					14'b01000100110010: oled_data = 16'b0111110101111011;
					14'b01011010110010: oled_data = 16'b1001010111111011;
					14'b01011100110010: oled_data = 16'b1100011011011101;
					14'b01100100110010: oled_data = 16'b1100111100011000;
					14'b01100110110010: oled_data = 16'b1001011000001110;
					14'b01101000110010: oled_data = 16'b1110011110011100;
					14'b01101010110010: oled_data = 16'b1110011110011100;
					14'b01101100110010: oled_data = 16'b1110011110011100;
					14'b01101110110010: oled_data = 16'b1110011110011100;
					14'b01110000110010: oled_data = 16'b1110011110011100;
					14'b01110010110010: oled_data = 16'b1110011110011100;
					14'b01110100110010: oled_data = 16'b1110011110011100;
					14'b01110110110010: oled_data = 16'b1110011110011100;
					14'b01111000110010: oled_data = 16'b1001011000001110;
					14'b01111010110010: oled_data = 16'b1100111100111000;
					14'b01000010110011: oled_data = 16'b1110011101111110;
					14'b01000100110011: oled_data = 16'b0110110100111010;
					14'b01000110110011: oled_data = 16'b1010111001111100;
					14'b01001000110011: oled_data = 16'b1011011001111100;
					14'b01001010110011: oled_data = 16'b1011011001111100;
					14'b01001100110011: oled_data = 16'b1011011001111100;
					14'b01001110110011: oled_data = 16'b1011011010011100;
					14'b01010000110011: oled_data = 16'b1011011010011100;
					14'b01010010110011: oled_data = 16'b1011011010011100;
					14'b01010100110011: oled_data = 16'b1011011001111100;
					14'b01010110110011: oled_data = 16'b1011011001111100;
					14'b01011000110011: oled_data = 16'b1011011001111100;
					14'b01011010110011: oled_data = 16'b0111010101011010;
					14'b01011100110011: oled_data = 16'b1100011011011101;
					14'b01100100110011: oled_data = 16'b1101111101111010;
					14'b01100110110011: oled_data = 16'b1000110111101101;
					14'b01101000110011: oled_data = 16'b1001011000001110;
					14'b01101010110011: oled_data = 16'b1001011000001110;
					14'b01101100110011: oled_data = 16'b1001011000001110;
					14'b01101110110011: oled_data = 16'b1000110111101110;
					14'b01110000110011: oled_data = 16'b1000110111101110;
					14'b01110010110011: oled_data = 16'b1001011000001110;
					14'b01110100110011: oled_data = 16'b1001011000001110;
					14'b01110110110011: oled_data = 16'b1001011000001110;
					14'b01111000110011: oled_data = 16'b1000110111101101;
					14'b01111010110011: oled_data = 16'b1101111101111010;
					14'b01000010110100: oled_data = 16'b1111011111011110;
					14'b01000100110100: oled_data = 16'b1011011010011100;
					14'b01000110110100: oled_data = 16'b1001111000111100;
					14'b01001000110100: oled_data = 16'b1010011000111100;
					14'b01001010110100: oled_data = 16'b1010011001011100;
					14'b01001100110100: oled_data = 16'b1001111000011100;
					14'b01001110110100: oled_data = 16'b0101010010111001;
					14'b01010000110100: oled_data = 16'b0100110010011001;
					14'b01010010110100: oled_data = 16'b1000110110111011;
					14'b01010100110100: oled_data = 16'b1010011001011100;
					14'b01010110110100: oled_data = 16'b1010011000111100;
					14'b01011000110100: oled_data = 16'b1010011000111100;
					14'b01011010110100: oled_data = 16'b1010011001011100;
					14'b01011100110100: oled_data = 16'b1110111110011110;
					14'b01100000110100: oled_data = 16'b1110111110111101;
					14'b01100010110100: oled_data = 16'b1011011010010011;
					14'b01100100110100: oled_data = 16'b1010111010010010;
					14'b01100110110100: oled_data = 16'b1010111001110010;
					14'b01101000110100: oled_data = 16'b1010111001110010;
					14'b01101010110100: oled_data = 16'b1010111001110010;
					14'b01101100110100: oled_data = 16'b1010111001110010;
					14'b01101110110100: oled_data = 16'b1100111100010111;
					14'b01110000110100: oled_data = 16'b1100111100010111;
					14'b01110010110100: oled_data = 16'b1010111001110010;
					14'b01110100110100: oled_data = 16'b1010111001110010;
					14'b01110110110100: oled_data = 16'b1010111001110010;
					14'b01111000110100: oled_data = 16'b1010111001110010;
					14'b01111010110100: oled_data = 16'b1010111010010010;
					14'b01111100110100: oled_data = 16'b1011011010110011;
					14'b01111110110100: oled_data = 16'b1110111110111101;
					14'b01001010110101: oled_data = 16'b1100011011011101;
					14'b01001100110101: oled_data = 16'b1001010111111011;
					14'b01001110110101: oled_data = 16'b0101010010111001;
					14'b01010000110101: oled_data = 16'b0100110010111001;
					14'b01010010110101: oled_data = 16'b1000010110111011;
					14'b01010100110101: oled_data = 16'b1011011001111100;
					14'b01100000110101: oled_data = 16'b1111011111011110;
					14'b01100010110101: oled_data = 16'b1011111011010101;
					14'b01100100110101: oled_data = 16'b1011011010110100;
					14'b01100110110101: oled_data = 16'b1011011010110100;
					14'b01101000110101: oled_data = 16'b1011011010110100;
					14'b01101010110101: oled_data = 16'b1011011010110100;
					14'b01101100110101: oled_data = 16'b1011011010110100;
					14'b01101110110101: oled_data = 16'b1011111011010101;
					14'b01110000110101: oled_data = 16'b1011111011010101;
					14'b01110010110101: oled_data = 16'b1011011010110100;
					14'b01110100110101: oled_data = 16'b1011011010110100;
					14'b01110110110101: oled_data = 16'b1011011010110100;
					14'b01111000110101: oled_data = 16'b1011011010110100;
					14'b01111010110101: oled_data = 16'b1011011010110011;
					14'b01111100110101: oled_data = 16'b1011111011010101;
					14'b01111110110101: oled_data = 16'b1111011111011110;
					14'b01001010110110: oled_data = 16'b1100111100011101;
					14'b01001100110110: oled_data = 16'b1011011010011100;
					14'b01001110110110: oled_data = 16'b1011111010111101;
					14'b01010000110110: oled_data = 16'b1011111011011101;
					14'b01010010110110: oled_data = 16'b1011011010111100;
					14'b01010100110110: oled_data = 16'b1100011011011101;
					14'b01010110110110: oled_data = 16'b1111011111011111;
				endcase
			end
			else if (menu_state > 4'd5) begin
				case ({x, y})
					14'b01001110011001: oled_data = 16'b1111011101111101;
					14'b01010000011001: oled_data = 16'b1110001110001101;
					14'b01010010011001: oled_data = 16'b1110010001010001;
					14'b01010100011001: oled_data = 16'b1111011111011110;
					14'b01001110011010: oled_data = 16'b1110110101110101;
					14'b01010000011010: oled_data = 16'b1100100000000000;
					14'b01010010011010: oled_data = 16'b1100100000000000;
					14'b01010100011010: oled_data = 16'b1111011011011010;
					14'b01110100011010: oled_data = 16'b1111011111011110;
					14'b01110110011010: oled_data = 16'b1100111011011101;
					14'b01111000011010: oled_data = 16'b1100011010011100;
					14'b01111010011010: oled_data = 16'b1110111110011110;
					14'b01001110011011: oled_data = 16'b1111011101011100;
					14'b01010000011011: oled_data = 16'b1101101001101001;
					14'b01010010011011: oled_data = 16'b1110001110001101;
					14'b01010100011011: oled_data = 16'b1111011110111110;
					14'b01110100011011: oled_data = 16'b1111011110111110;
					14'b01110110011011: oled_data = 16'b0101001111111000;
					14'b01111000011011: oled_data = 16'b0011101101010111;
					14'b01111010011011: oled_data = 16'b1100111010111101;
					14'b01001010011100: oled_data = 16'b1111111111011110;
					14'b01001100011100: oled_data = 16'b1110110111110111;
					14'b01001110011100: oled_data = 16'b1101101100101100;
					14'b01010000011100: oled_data = 16'b1101000110100110;
					14'b01010010011100: oled_data = 16'b1110110110110110;
					14'b01110100011100: oled_data = 16'b1111011111011110;
					14'b01110110011100: oled_data = 16'b0101110000011000;
					14'b01111000011100: oled_data = 16'b0011101101110111;
					14'b01111010011100: oled_data = 16'b1100111011011101;
					14'b01001010011101: oled_data = 16'b1110001110001101;
					14'b01001100011101: oled_data = 16'b1100100000100000;
					14'b01001110011101: oled_data = 16'b1100100000000000;
					14'b01010000011101: oled_data = 16'b1100100000000000;
					14'b01010010011101: oled_data = 16'b1101000101100101;
					14'b01010100011101: oled_data = 16'b1111011110111110;
					14'b01110000011101: oled_data = 16'b1011111001011100;
					14'b01110010011101: oled_data = 16'b1001010110011011;
					14'b01110100011101: oled_data = 16'b1100011010111101;
					14'b01110110011101: oled_data = 16'b0101110000111000;
					14'b01111000011101: oled_data = 16'b0011101101110111;
					14'b01111010011101: oled_data = 16'b1100111011011101;
					14'b01001000011110: oled_data = 16'b1111011011111011;
					14'b01001010011110: oled_data = 16'b1100100001100001;
					14'b01001100011110: oled_data = 16'b1110010000110000;
					14'b01001110011110: oled_data = 16'b1101000010000010;
					14'b01010000011110: oled_data = 16'b1100100000000000;
					14'b01010010011110: oled_data = 16'b1100100000000000;
					14'b01010100011110: oled_data = 16'b1110110100010011;
					14'b01110000011110: oled_data = 16'b0111010011011001;
					14'b01110010011110: oled_data = 16'b0010101100010111;
					14'b01110100011110: oled_data = 16'b1001110110011011;
					14'b01110110011110: oled_data = 16'b0110010001011001;
					14'b01111000011110: oled_data = 16'b0011101101110111;
					14'b01111010011110: oled_data = 16'b1100111011011101;
					14'b01001000011111: oled_data = 16'b1110110101010100;
					14'b01001010011111: oled_data = 16'b1101000110100110;
					14'b01001100011111: oled_data = 16'b1110110110010101;
					14'b01001110011111: oled_data = 16'b1100100000000000;
					14'b01010000011111: oled_data = 16'b1101000011000011;
					14'b01010010011111: oled_data = 16'b1101101010101010;
					14'b01010100011111: oled_data = 16'b1100100001000001;
					14'b01010110011111: oled_data = 16'b1101000110000110;
					14'b01011000011111: oled_data = 16'b1110111000011000;
					14'b01110000011111: oled_data = 16'b0111110011111010;
					14'b01110010011111: oled_data = 16'b0011001100110111;
					14'b01110100011111: oled_data = 16'b1001110110111011;
					14'b01110110011111: oled_data = 16'b0110010001011001;
					14'b01111000011111: oled_data = 16'b0011101101110111;
					14'b01111010011111: oled_data = 16'b1100111011011101;
					14'b01001000100000: oled_data = 16'b1111011110011101;
					14'b01001010100000: oled_data = 16'b1111011101011100;
					14'b01001100100000: oled_data = 16'b1110010001010000;
					14'b01001110100000: oled_data = 16'b1100100000000000;
					14'b01010000100000: oled_data = 16'b1101000111000111;
					14'b01010100100000: oled_data = 16'b1110111000111000;
					14'b01010110100000: oled_data = 16'b1110001111001110;
					14'b01011000100000: oled_data = 16'b1110111001011000;
					14'b01101010100000: oled_data = 16'b1011111001111100;
					14'b01101100100000: oled_data = 16'b0110110010011001;
					14'b01101110100000: oled_data = 16'b1010010111011011;
					14'b01110000100000: oled_data = 16'b0111110011111010;
					14'b01110010100000: oled_data = 16'b0011001100110111;
					14'b01110100100000: oled_data = 16'b1001110110111011;
					14'b01110110100000: oled_data = 16'b0110010001011001;
					14'b01111000100000: oled_data = 16'b0011101101110111;
					14'b01111010100000: oled_data = 16'b1100111011011101;
					14'b01001100100001: oled_data = 16'b1101101010001010;
					14'b01001110100001: oled_data = 16'b1100100010000010;
					14'b01010000100001: oled_data = 16'b1100100001100001;
					14'b01010010100001: oled_data = 16'b1110010010010001;
					14'b01101010100001: oled_data = 16'b1001110110111011;
					14'b01101100100001: oled_data = 16'b0010101100010111;
					14'b01101110100001: oled_data = 16'b0111110011111010;
					14'b01110000100001: oled_data = 16'b0111110100011010;
					14'b01110010100001: oled_data = 16'b0011001100110111;
					14'b01110100100001: oled_data = 16'b1001110110111011;
					14'b01110110100001: oled_data = 16'b0110010001011001;
					14'b01111000100001: oled_data = 16'b0011101101110111;
					14'b01111010100001: oled_data = 16'b1100111011011101;
					14'b01001010100010: oled_data = 16'b1111111111011110;
					14'b01001100100010: oled_data = 16'b1101000011100011;
					14'b01001110100010: oled_data = 16'b1110010010110010;
					14'b01010000100010: oled_data = 16'b1110010011010010;
					14'b01010010100010: oled_data = 16'b1100100000100000;
					14'b01010100100010: oled_data = 16'b1110110100010011;
					14'b01100100100010: oled_data = 16'b1111011111011110;
					14'b01100110100010: oled_data = 16'b1110111110111110;
					14'b01101000100010: oled_data = 16'b1111011110111110;
					14'b01101010100010: oled_data = 16'b1010010111011011;
					14'b01101100100010: oled_data = 16'b0011001100110111;
					14'b01101110100010: oled_data = 16'b1000010100011010;
					14'b01110000100010: oled_data = 16'b0111110100011010;
					14'b01110010100010: oled_data = 16'b0011001100110111;
					14'b01110100100010: oled_data = 16'b1001110110111011;
					14'b01110110100010: oled_data = 16'b0110010001011001;
					14'b01111000100010: oled_data = 16'b0011101101110111;
					14'b01111010100010: oled_data = 16'b1100111011011101;
					14'b01001010100011: oled_data = 16'b1110010011110011;
					14'b01001100100011: oled_data = 16'b1100100000100000;
					14'b01001110100011: oled_data = 16'b1111011010111010;
					14'b01010010100011: oled_data = 16'b1101000101100101;
					14'b01010100100011: oled_data = 16'b1110010000110000;
					14'b01100100100011: oled_data = 16'b1100111011011101;
					14'b01100110100011: oled_data = 16'b0100101111011000;
					14'b01101000100011: oled_data = 16'b0111010010111001;
					14'b01101010100011: oled_data = 16'b1001110110111011;
					14'b01101100100011: oled_data = 16'b0011001100110111;
					14'b01101110100011: oled_data = 16'b1000010100011010;
					14'b01110000100011: oled_data = 16'b0111110100011010;
					14'b01110010100011: oled_data = 16'b0011001100110111;
					14'b01110100100011: oled_data = 16'b1001110110111011;
					14'b01110110100011: oled_data = 16'b0110010001011001;
					14'b01111000100011: oled_data = 16'b0011101101110111;
					14'b01111010100011: oled_data = 16'b1100111011011101;
					14'b01001000100100: oled_data = 16'b1110111000010111;
					14'b01001010100100: oled_data = 16'b1100100000100000;
					14'b01001100100100: oled_data = 16'b1110010001110001;
					14'b01010010100100: oled_data = 16'b1101000101100101;
					14'b01010100100100: oled_data = 16'b1110010001010000;
					14'b01100100100100: oled_data = 16'b1100011010111101;
					14'b01100110100100: oled_data = 16'b0011001101010111;
					14'b01101000100100: oled_data = 16'b0110010000111001;
					14'b01101010100100: oled_data = 16'b1001110110111011;
					14'b01101100100100: oled_data = 16'b0011001100110111;
					14'b01101110100100: oled_data = 16'b1000010100011010;
					14'b01110000100100: oled_data = 16'b0111110100011010;
					14'b01110010100100: oled_data = 16'b0011001100110111;
					14'b01110100100100: oled_data = 16'b1001110110111011;
					14'b01110110100100: oled_data = 16'b0110010000111001;
					14'b01111000100100: oled_data = 16'b0011101101010111;
					14'b01111010100100: oled_data = 16'b1100111011011101;
					14'b01000110100101: oled_data = 16'b1111011100011011;
					14'b01001000100101: oled_data = 16'b1101000010100010;
					14'b01001010100101: oled_data = 16'b1101101100001100;
					14'b01010010100101: oled_data = 16'b1101000100100100;
					14'b01010100100101: oled_data = 16'b1110010000110000;
					14'b01100100100101: oled_data = 16'b1110111110011110;
					14'b01100110100101: oled_data = 16'b1100111011011101;
					14'b01101000100101: oled_data = 16'b1101011100011101;
					14'b01101010100101: oled_data = 16'b1110011101011110;
					14'b01101100100101: oled_data = 16'b1100111011011101;
					14'b01101110100101: oled_data = 16'b1101111100111110;
					14'b01110000100101: oled_data = 16'b1101111100111101;
					14'b01110010100101: oled_data = 16'b1100111011011101;
					14'b01110100100101: oled_data = 16'b1110011101111110;
					14'b01110110100101: oled_data = 16'b1101011100011101;
					14'b01111000100101: oled_data = 16'b1100111011011101;
					14'b01111010100101: oled_data = 16'b1110111110111110;
					14'b01000110100110: oled_data = 16'b1111011100011011;
					14'b01001000100110: oled_data = 16'b1110010000001111;
					14'b01001010100110: oled_data = 16'b1111011110111110;
					14'b01010010100110: oled_data = 16'b1110010011010010;
					14'b01010100100110: oled_data = 16'b1110111001011000;
					14'b01000100101010: oled_data = 16'b1110111100111011;
					14'b01000110101010: oled_data = 16'b1100110111010100;
					14'b01000010101011: oled_data = 16'b1111011111011110;
					14'b01000100101011: oled_data = 16'b1010001110101010;
					14'b01000110101011: oled_data = 16'b0111100101100000;
					14'b01001000101011: oled_data = 16'b1100010101010010;
					14'b01101110101011: oled_data = 16'b1111111110111110;
					14'b01110000101011: oled_data = 16'b1111111110111110;
					14'b01000100101100: oled_data = 16'b1101111001110111;
					14'b01000110101100: oled_data = 16'b1000101001000011;
					14'b01001000101100: oled_data = 16'b0111100110000000;
					14'b01001010101100: oled_data = 16'b1100110101110011;
					14'b01101010101100: oled_data = 16'b1111111111011110;
					14'b01101100101100: oled_data = 16'b1111111000111011;
					14'b01101110101100: oled_data = 16'b1111110011111001;
					14'b01110000101100: oled_data = 16'b1111110100011001;
					14'b01110010101100: oled_data = 16'b1111111000111011;
					14'b01110100101100: oled_data = 16'b1111111111011110;
					14'b01000110101101: oled_data = 16'b1110011010111001;
					14'b01001000101101: oled_data = 16'b1000101001100100;
					14'b01001010101101: oled_data = 16'b0111100110100000;
					14'b01001100101101: oled_data = 16'b1100110110110100;
					14'b01101010101101: oled_data = 16'b1111111001111100;
					14'b01101100101101: oled_data = 16'b1111110001111000;
					14'b01101110101101: oled_data = 16'b1111110011111001;
					14'b01110000101101: oled_data = 16'b1111110010111000;
					14'b01110010101101: oled_data = 16'b1111110001111000;
					14'b01110100101101: oled_data = 16'b1111111001111100;
					14'b01001000101110: oled_data = 16'b1110011011011010;
					14'b01001010101110: oled_data = 16'b1000101010000101;
					14'b01001100101110: oled_data = 16'b0111100110100000;
					14'b01001110101110: oled_data = 16'b1101010111110101;
					14'b01101010101110: oled_data = 16'b1111110101111010;
					14'b01101100101110: oled_data = 16'b1111110100111001;
					14'b01101110101110: oled_data = 16'b1111111000011011;
					14'b01110000101110: oled_data = 16'b1111110110011010;
					14'b01110010101110: oled_data = 16'b1111110100111001;
					14'b01110100101110: oled_data = 16'b1111110101111010;
					14'b01001010101111: oled_data = 16'b1110011100011010;
					14'b01001100101111: oled_data = 16'b1001001010100101;
					14'b01001110101111: oled_data = 16'b0111100111000001;
					14'b01010000101111: oled_data = 16'b1101011000010110;
					14'b01101010101111: oled_data = 16'b1111110110111010;
					14'b01101100101111: oled_data = 16'b1111110110111010;
					14'b01101110101111: oled_data = 16'b1111110011011000;
					14'b01110000101111: oled_data = 16'b1111110100011001;
					14'b01110010101111: oled_data = 16'b1111110111011010;
					14'b01110100101111: oled_data = 16'b1111110110111010;
					14'b01001100110000: oled_data = 16'b1110111100111011;
					14'b01001110110000: oled_data = 16'b1001001011000110;
					14'b01010000110000: oled_data = 16'b1000000111100001;
					14'b01010010110000: oled_data = 16'b1101111001110111;
					14'b01010100110000: oled_data = 16'b1110111101011100;
					14'b01010110110000: oled_data = 16'b1010001101101001;
					14'b01011000110000: oled_data = 16'b1011110011001111;
					14'b01101010110000: oled_data = 16'b1111111000011011;
					14'b01101100110000: oled_data = 16'b1111110110011010;
					14'b01101110110000: oled_data = 16'b1111110010011000;
					14'b01110000110000: oled_data = 16'b1111110010011000;
					14'b01110010110000: oled_data = 16'b1111110110111010;
					14'b01110100110000: oled_data = 16'b1111111000011011;
					14'b01001110110001: oled_data = 16'b1110111101011100;
					14'b01010000110001: oled_data = 16'b1001101100000111;
					14'b01010010110001: oled_data = 16'b1000101001000011;
					14'b01010100110001: oled_data = 16'b1001001011000101;
					14'b01010110110001: oled_data = 16'b0111100110000000;
					14'b01011000110001: oled_data = 16'b0111100110100000;
					14'b01011010110001: oled_data = 16'b1011110011001111;
					14'b01011100110001: oled_data = 16'b1111011111011110;
					14'b01101000110001: oled_data = 16'b1111111111011110;
					14'b01101010110001: oled_data = 16'b1111110111011010;
					14'b01101100110001: oled_data = 16'b1111111011011100;
					14'b01101110110001: oled_data = 16'b1111111010011100;
					14'b01110000110001: oled_data = 16'b1111111010011100;
					14'b01110010110001: oled_data = 16'b1111111011011100;
					14'b01110100110001: oled_data = 16'b1111110111011010;
					14'b01110110110001: oled_data = 16'b1111111111011110;
					14'b01010000110010: oled_data = 16'b1110011010111001;
					14'b01010010110010: oled_data = 16'b1000000111100001;
					14'b01010100110010: oled_data = 16'b0111100110100000;
					14'b01010110110010: oled_data = 16'b1000000111000001;
					14'b01011000110010: oled_data = 16'b0111100110100000;
					14'b01011010110010: oled_data = 16'b1000101001000011;
					14'b01011100110010: oled_data = 16'b1110111101011100;
					14'b01101000110010: oled_data = 16'b1111111110011110;
					14'b01101010110010: oled_data = 16'b1111110110011010;
					14'b01101100110010: oled_data = 16'b1111111010011100;
					14'b01101110110010: oled_data = 16'b1111111000011011;
					14'b01110000110010: oled_data = 16'b1111111000011011;
					14'b01110010110010: oled_data = 16'b1111111010011100;
					14'b01110100110010: oled_data = 16'b1111110110011010;
					14'b01110110110010: oled_data = 16'b1111111110011110;
					14'b01001110110011: oled_data = 16'b1110111101111100;
					14'b01010000110011: oled_data = 16'b1001101100101000;
					14'b01010010110011: oled_data = 16'b0111100110100000;
					14'b01010100110011: oled_data = 16'b1000000111000001;
					14'b01010110110011: oled_data = 16'b0111100111000000;
					14'b01011000110011: oled_data = 16'b1000000111100001;
					14'b01011010110011: oled_data = 16'b1101011000010110;
					14'b01100110110011: oled_data = 16'b1111111111011111;
					14'b01101000110011: oled_data = 16'b1111111001011011;
					14'b01101010110011: oled_data = 16'b1111110011011000;
					14'b01101100110011: oled_data = 16'b1111111010111100;
					14'b01101110110011: oled_data = 16'b1111111010011100;
					14'b01110000110011: oled_data = 16'b1111111010011100;
					14'b01110010110011: oled_data = 16'b1111111010111100;
					14'b01110100110011: oled_data = 16'b1111110011011000;
					14'b01110110110011: oled_data = 16'b1111111001011011;
					14'b01111000110011: oled_data = 16'b1111111111011111;
					14'b01001110110100: oled_data = 16'b1110011010111001;
					14'b01010000110100: oled_data = 16'b1000001000000010;
					14'b01010010110100: oled_data = 16'b0111100111000001;
					14'b01010100110100: oled_data = 16'b0111100111000000;
					14'b01010110110100: oled_data = 16'b1000001000000010;
					14'b01011000110100: oled_data = 16'b1101010111010101;
					14'b01100110110100: oled_data = 16'b1111111110111110;
					14'b01101000110100: oled_data = 16'b1111110011111001;
					14'b01101010110100: oled_data = 16'b1111110010111000;
					14'b01101100110100: oled_data = 16'b1111110011011000;
					14'b01101110110100: oled_data = 16'b1111110100111001;
					14'b01110000110100: oled_data = 16'b1111110100111001;
					14'b01110010110100: oled_data = 16'b1111110011011000;
					14'b01110100110100: oled_data = 16'b1111110010111000;
					14'b01110110110100: oled_data = 16'b1111110011111001;
					14'b01111000110100: oled_data = 16'b1111111110111110;
					14'b01001000110101: oled_data = 16'b1111011111011110;
					14'b01001010110101: oled_data = 16'b1110011011111010;
					14'b01001100110101: oled_data = 16'b1100010101010010;
					14'b01001110110101: oled_data = 16'b1100110110010011;
					14'b01010000110101: oled_data = 16'b1011010001101110;
					14'b01010010110101: oled_data = 16'b1000000111100001;
					14'b01010100110101: oled_data = 16'b1000001000000010;
					14'b01010110110101: oled_data = 16'b1010001111001010;
					14'b01011000110101: oled_data = 16'b1101010111110101;
					14'b01011010110101: oled_data = 16'b1101111010011000;
					14'b01011100110101: oled_data = 16'b1111011111011110;
					14'b01100110110101: oled_data = 16'b1111111110011110;
					14'b01101000110101: oled_data = 16'b1111110011111001;
					14'b01101010110101: oled_data = 16'b1111110010011000;
					14'b01101100110101: oled_data = 16'b1111110010011000;
					14'b01101110110101: oled_data = 16'b1111110100111001;
					14'b01110000110101: oled_data = 16'b1111110100111001;
					14'b01110010110101: oled_data = 16'b1111110010011000;
					14'b01110100110101: oled_data = 16'b1111110010011000;
					14'b01110110110101: oled_data = 16'b1111110011111001;
					14'b01111000110101: oled_data = 16'b1111111110011110;
					14'b01001000110110: oled_data = 16'b1111011101111101;
					14'b01001010110110: oled_data = 16'b1101111001010111;
					14'b01001100110110: oled_data = 16'b1110011010111001;
					14'b01001110110110: oled_data = 16'b1111011110011101;
					14'b01010000110110: oled_data = 16'b1100110110010011;
					14'b01010010110110: oled_data = 16'b1001101101001000;
					14'b01010100110110: oled_data = 16'b1101010111110101;
					14'b01010110110110: oled_data = 16'b1101011000010110;
					14'b01011000110110: oled_data = 16'b1101111001110111;
					14'b01011010110110: oled_data = 16'b1111011101111101;
					14'b01011100110110: oled_data = 16'b1111011111011110;
					14'b01100110110110: oled_data = 16'b1111111111011110;
					14'b01101000110110: oled_data = 16'b1111111011011100;
					14'b01101010110110: oled_data = 16'b1111111010111100;
					14'b01101100110110: oled_data = 16'b1111111010111100;
					14'b01101110110110: oled_data = 16'b1111111011111101;
					14'b01110000110110: oled_data = 16'b1111111011111101;
					14'b01110010110110: oled_data = 16'b1111111010111100;
					14'b01110100110110: oled_data = 16'b1111111010111100;
					14'b01110110110110: oled_data = 16'b1111111011011100;
					14'b01111000110110: oled_data = 16'b1111111111011110;
					14'b01001110110111: oled_data = 16'b1110111101111100;
					14'b01010000110111: oled_data = 16'b1101111010011000;
					14'b01010010110111: oled_data = 16'b1101111001010111;
					14'b01010100110111: oled_data = 16'b1111011110111110;
					14'b01010110110111: oled_data = 16'b1111011110111110;
				endcase
			end
		end
	end

endmodule