`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/25/2023 05:03:22 PM
// Design Name: 
// Module Name: audio_game_oled
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module audio_game_oled(
    input clock, clk_os, clk_display, clk_pos, btnC, btnU,
    input [10:0] num, 
    input [6:0] x,y,
    output [15:0] oled_data
    );
    
    parameter reg gravity = 5;
    reg flag = 0;
    reg [4:0] y_acc;
    wire [4:0] y_acceleration;
    wire x_move;
    wire [31:0] offset;
    wire [1:0] stop_x;
    always @ (posedge clock) begin
        if (num >= 0 && num < 205)
            begin  
                y_acc <= 0;
                flag <= 0;
            end
        else if (num >= 205 && num < 409)
            begin
                y_acc <= 50;
                flag <= 1;
            end
        else if (num >= 409 && num < 614)
            begin
                y_acc <= 45;
                flag <= 1;            
            end
        else if (num >= 614 && num < 819)
            begin
                y_acc <= 40;
                flag <= 1;            
            end
        else if (num >= 819 && num < 1024)
            begin 
                y_acc <= 35;
                flag <= 1;            
            end
        else if (num >= 1024 && num < 1229)
            begin 
                y_acc <= 30;
                flag <= 1;            
            end
        else if (num >= 1229 && num < 1434)
            begin
                y_acc <= 25;
                flag <= 1;            
            end
        else if (num >= 1434 && num < 1638)
            begin
                y_acc <= 20;
                flag <= 1;            
            end
        else if (num >= 1638 && num < 1842)
            begin
                y_acc <= 15;
                flag <= 1;            
            end
        else if (num >= 1842 && num <= 2047)
            begin 
                y_acc <= 10;
                flag <= 1;            
            end
    end
    
    assign y_acceleration = y_acc;
    assign x_move = flag && stop_x;
    
    check_x_offset x_offset(clk_os, x_move, btnC, offset);
    output_display oled(clk_display, clk_pos, btnC, btnU, y_acceleration, x,y,offset, stop_x, oled_data);
endmodule


module check_x_offset(
    input clk_os, x_move, btnC,
    output reg [31:0] offset = 0
);

    parameter max_offset = 1406;
    always @ (posedge clk_os) begin
        if (x_move) begin
            offset <= (offset == max_offset) || btnC ? 0 : offset + 1;
        end
        
        else offset <= btnC ? 0 : offset;
    end
    
endmodule

module output_display(
    input clk_display, clk_pos, btnC, btnU,
    input [4:0] y_acc,
    input [6:0] x,y,
    input [31:0] offset,
    output reg [1:0] stop_x = 1,
    output reg [15:0] oled_data
);

    wire [15:0] data [0:15019];
    wire [31:0] index;
    assign index = (x * 10) + (y - 54) + (10 * offset);
    
    parameter square_size = 3;
    parameter max_y_pos = 3;
    parameter min_y_pos = 60;
    
    wire square_pos;
    //initial position of ball
    reg [6:0] x_pos = 25;
    reg [6:0] y_pos = 20; 
    
    reg [31:0] count = 0;
    
    // boolean logics 
    wire hit_top, hit_bottom, hit_right, on_land;
    wire index_to_check_right;
    wire [31:0] index_to_check_bottom [0:6];
    wire [31:0] col_num [0:29];
    //death screen
    wire [15:0] death_oled;
    
    //score screen
    wire [15:0] score_oled;
    reg score_flag = 0;
    
    //score system
    reg [4:0] prev_blk;
    reg [4:0] curr_blk;
    reg [4:0] score = 0;
    
    //assign all boolean logic here
    assign hit_top = (y_pos <= max_y_pos);
    assign hit_bottom = (y_pos >= min_y_pos);
    assign index_to_check_right = 290 + (y_pos + square_size - 54) + 10 * offset;
    assign index_to_check_bottom[0] = 220 + offset * 10;
    assign index_to_check_bottom[1] = 230 + offset * 10;
    assign index_to_check_bottom[2] = 240 + offset * 10;
    assign index_to_check_bottom[3] = 250 + offset * 10;
    assign index_to_check_bottom[4] = 260 + offset * 10;
    assign index_to_check_bottom[5] = 270 + offset * 10;
    assign index_to_check_bottom[6] = 280 + offset * 10;
    assign hit_right = (y_pos > 50) && (data[index_to_check_right] == 16'b0);
    assign on_land = (y_pos == 50) && (data[index_to_check_bottom[0]] == 16'b0 || 
                                       data[index_to_check_bottom[1]] == 16'b0 || 
                                       data[index_to_check_bottom[2]] == 16'b0 || 
                                       data[index_to_check_bottom[3]] == 16'b0 || 
                                       data[index_to_check_bottom[4]] == 16'b0 || 
                                       data[index_to_check_bottom[5]] == 16'b0 || 
                                       data[index_to_check_bottom[6]] == 16'b0);
    assign col_num[0] = offset <= 7;
    assign col_num[1] = (offset >= 40 - 28) && (offset <= 72 - 22);
    assign col_num[2] = (offset >= 93 - 28) && (offset <= 121 - 22);
    assign col_num[3] = (offset >= 141 - 28) && (offset <= 178 - 22);
    assign col_num[4] = (offset >= 202 - 28) && (offset <= 221 - 22);
    assign col_num[5] = (offset >= 232 - 28) && (offset <= 252 - 22);
    assign col_num[6] = (offset >= 270 - 28) && (offset <= 302 - 22);
    assign col_num[7] = (offset >= 327 - 28) && (offset <= 362 - 22);
    assign col_num[8] = (offset >= 379 - 28) && (offset <= 416 - 22);
    assign col_num[9] = (offset >= 427 - 28) && (offset <= 466 - 22);
    assign col_num[10] = (offset >= 480 - 28) && (offset <= 505 - 22);
    assign col_num[11] = (offset >= 523 - 28) && (offset <= 562 - 22);
    assign col_num[12] = (offset >= 580 - 28) && (offset <= 617 - 22);
    assign col_num[13] = (offset >= 628 - 28) && (offset <= 667 - 22);
    assign col_num[14] = (offset >= 685 - 28) && (offset <= 709 - 22);
    assign col_num[15] = (offset >= 722 - 28) && (offset <= 741 - 22);
    assign col_num[16] = (offset >= 755 - 28) && (offset <= 787 - 22);
    assign col_num[17] = (offset >= 813 - 28) && (offset <= 832 - 22);
    assign col_num[18] = (offset >= 847 - 28) && (offset <= 870 - 22);
    assign col_num[19] = (offset >= 886 - 28) && (offset <= 923 - 22);
    assign col_num[20] = (offset >= 949 - 28) && (offset <= 985 - 22);
    assign col_num[21] = (offset >= 1007 - 28) && (offset <= 1036 - 22);
    assign col_num[22] = (offset >= 1061 - 28) && (offset <= 1086 - 22);
    assign col_num[23] = (offset >= 1107 - 28) && (offset <= 1128 - 22);
    assign col_num[24] = (offset >= 1143 - 28) && (offset <= 1182 - 22);
    assign col_num[25] = (offset >= 1196 - 28) && (offset <= 1225 - 22);
    assign col_num[26] = (offset >= 1240 - 28) && (offset <= 1278 - 22);
    assign col_num[27] = (offset >= 1298 - 28) && (offset <= 1329 - 22);
    assign col_num[28] = (offset >= 1341 - 28) && (offset <= 1379 - 22);
    assign col_num[29] = (offset >= 1390 - 28) && (offset <= 1428 - 22);
    
    
    
    
    //output logic of x,y coordinates to render the square
    assign square_pos  = (x >= x_pos - square_size && x <= x_pos + square_size) &&
                         (y >= y_pos - square_size && y <= y_pos + square_size);
                         
                        
    always @(posedge clk_display) begin
        stop_x <= hit_right || hit_bottom ? 0 : 1;
        oled_data <= score_flag ? score_oled : hit_bottom ? death_oled : square_pos ? 16'b0 : y > 53 ? data[index] : ~16'b0;
    end
    
    always @(posedge clk_pos) begin
        score_flag <= btnC ? 0 : btnU ? 1 : score_flag;
        if (y_acc > 0) begin
            count <= count >= y_acc - 1 ? 0 : count + 1;
            y_pos <= btnC ? 20 : (count == y_acc - 1? (hit_top ? max_y_pos : hit_bottom ? min_y_pos : y_pos - 1) : y_pos);
        end
        
        else begin
            count <= count >= 14 ? 0 : count + 1;
            y_pos <= btnC ? 20 : (count == 14 ? (hit_bottom ? min_y_pos : on_land ? 50 : y_pos + 1) : y_pos);
        end
        if (btnC) begin
            score <= 0;
            prev_blk <= 1;
            curr_blk <= 1;
        end
        
        else begin
            if(on_land) begin
            curr_blk <= col_num[0] ? 1 :
                       col_num[1] ? 2 :
                       col_num[2] ? 3 :
                       col_num[3] ? 4 :
                       col_num[4] ? 5 :
                       col_num[5] ? 6 :
                       col_num[6] ? 7 :
                       col_num[7] ? 8 :
                       col_num[8] ? 9 :
                       col_num[9] ? 10 :
                       col_num[10] ? 11 :
                       col_num[11] ? 12 :
                       col_num[12] ? 13 :
                       col_num[13] ? 14 :
                       col_num[14] ? 15 :
                       col_num[15] ? 16 :
                       col_num[16] ? 17 :
                       col_num[17] ? 18 :
                       col_num[18] ? 19 :
                       col_num[19] ? 20 :
                       col_num[20] ? 21 :
                       col_num[21] ? 22 :
                       col_num[22] ? 23 :
                       col_num[23] ? 24 :
                       col_num[24] ? 25 :
                       col_num[25] ? 26 :
                       col_num[26] ? 27 :
                       col_num[27] ? 28 :
                       col_num[28] ? 29 :
                       col_num[29] ? 30 : 0;
            score <= curr_blk != prev_blk ? score + 1 : score;
            prev_blk <= curr_blk;
            end   
        end           
    end
    
    
    death_image d1(.x(x), .y(y), .oled_data(death_oled));
    oled_score score_display(clk_display, score,x,y,score_oled );
    assign data[0] = 16'b0;
    assign data[1] = 16'b0;
    assign data[2] = 16'b0;
    assign data[3] = 16'b0;
    assign data[4] = 16'b0;
    assign data[5] = 16'b0;
    assign data[6] = 16'b0;
    assign data[7] = 16'b0;
    assign data[8] = 16'b0;
    assign data[9] = 16'b0;
    assign data[10] = 16'b0;
    assign data[11] = 16'b0;
    assign data[12] = 16'b0;
    assign data[13] = 16'b0;
    assign data[14] = 16'b0;
    assign data[15] = 16'b0;
    assign data[16] = 16'b0;
    assign data[17] = 16'b0;
    assign data[18] = 16'b0;
    assign data[19] = 16'b0;
    assign data[20] = 16'b0;
    assign data[21] = 16'b0;
    assign data[22] = ~16'b0;
    assign data[23] = ~16'b0;
    assign data[24] = ~16'b0;
    assign data[25] = ~16'b0;
    assign data[26] = ~16'b0;
    assign data[27] = ~16'b0;
    assign data[28] = ~16'b0;
    assign data[29] = ~16'b0;
    assign data[30] = 16'b0;
    assign data[31] = 16'b0;
    assign data[32] = ~16'b0;
    assign data[33] = ~16'b0;
    assign data[34] = ~16'b0;
    assign data[35] = ~16'b0;
    assign data[36] = ~16'b0;
    assign data[37] = ~16'b0;
    assign data[38] = ~16'b0;
    assign data[39] = ~16'b0;
    assign data[40] = 16'b0;
    assign data[41] = 16'b0;
    assign data[42] = ~16'b0;
    assign data[43] = ~16'b0;
    assign data[44] = ~16'b0;
    assign data[45] = ~16'b0;
    assign data[46] = ~16'b0;
    assign data[47] = ~16'b0;
    assign data[48] = ~16'b0;
    assign data[49] = ~16'b0;
    assign data[50] = 16'b0;
    assign data[51] = 16'b0;
    assign data[52] = ~16'b0;
    assign data[53] = ~16'b0;
    assign data[54] = ~16'b0;
    assign data[55] = ~16'b0;
    assign data[56] = ~16'b0;
    assign data[57] = ~16'b0;
    assign data[58] = ~16'b0;
    assign data[59] = ~16'b0;
    assign data[60] = 16'b0;
    assign data[61] = 16'b0;
    assign data[62] = ~16'b0;
    assign data[63] = ~16'b0;
    assign data[64] = ~16'b0;
    assign data[65] = ~16'b0;
    assign data[66] = ~16'b0;
    assign data[67] = ~16'b0;
    assign data[68] = ~16'b0;
    assign data[69] = ~16'b0;
    assign data[70] = 16'b0;
    assign data[71] = 16'b0;
    assign data[72] = ~16'b0;
    assign data[73] = ~16'b0;
    assign data[74] = ~16'b0;
    assign data[75] = ~16'b0;
    assign data[76] = ~16'b0;
    assign data[77] = ~16'b0;
    assign data[78] = ~16'b0;
    assign data[79] = ~16'b0;
    assign data[80] = 16'b0;
    assign data[81] = 16'b0;
    assign data[82] = ~16'b0;
    assign data[83] = ~16'b0;
    assign data[84] = ~16'b0;
    assign data[85] = ~16'b0;
    assign data[86] = ~16'b0;
    assign data[87] = ~16'b0;
    assign data[88] = ~16'b0;
    assign data[89] = ~16'b0;
    assign data[90] = 16'b0;
    assign data[91] = 16'b0;
    assign data[92] = ~16'b0;
    assign data[93] = ~16'b0;
    assign data[94] = ~16'b0;
    assign data[95] = ~16'b0;
    assign data[96] = ~16'b0;
    assign data[97] = ~16'b0;
    assign data[98] = ~16'b0;
    assign data[99] = ~16'b0;
    assign data[100] = 16'b0;
    assign data[101] = 16'b0;
    assign data[102] = ~16'b0;
    assign data[103] = ~16'b0;
    assign data[104] = ~16'b0;
    assign data[105] = ~16'b0;
    assign data[106] = ~16'b0;
    assign data[107] = ~16'b0;
    assign data[108] = ~16'b0;
    assign data[109] = ~16'b0;
    assign data[110] = 16'b0;
    assign data[111] = 16'b0;
    assign data[112] = ~16'b0;
    assign data[113] = ~16'b0;
    assign data[114] = ~16'b0;
    assign data[115] = ~16'b0;
    assign data[116] = ~16'b0;
    assign data[117] = ~16'b0;
    assign data[118] = ~16'b0;
    assign data[119] = ~16'b0;
    assign data[120] = 16'b0;
    assign data[121] = 16'b0;
    assign data[122] = ~16'b0;
    assign data[123] = ~16'b0;
    assign data[124] = ~16'b0;
    assign data[125] = ~16'b0;
    assign data[126] = ~16'b0;
    assign data[127] = ~16'b0;
    assign data[128] = ~16'b0;
    assign data[129] = ~16'b0;
    assign data[130] = 16'b0;
    assign data[131] = 16'b0;
    assign data[132] = ~16'b0;
    assign data[133] = ~16'b0;
    assign data[134] = ~16'b0;
    assign data[135] = ~16'b0;
    assign data[136] = ~16'b0;
    assign data[137] = ~16'b0;
    assign data[138] = ~16'b0;
    assign data[139] = ~16'b0;
    assign data[140] = 16'b0;
    assign data[141] = 16'b0;
    assign data[142] = ~16'b0;
    assign data[143] = ~16'b0;
    assign data[144] = ~16'b0;
    assign data[145] = ~16'b0;
    assign data[146] = ~16'b0;
    assign data[147] = ~16'b0;
    assign data[148] = ~16'b0;
    assign data[149] = ~16'b0;
    assign data[150] = 16'b0;
    assign data[151] = 16'b0;
    assign data[152] = ~16'b0;
    assign data[153] = ~16'b0;
    assign data[154] = ~16'b0;
    assign data[155] = ~16'b0;
    assign data[156] = ~16'b0;
    assign data[157] = ~16'b0;
    assign data[158] = ~16'b0;
    assign data[159] = ~16'b0;
    assign data[160] = 16'b0;
    assign data[161] = 16'b0;
    assign data[162] = ~16'b0;
    assign data[163] = ~16'b0;
    assign data[164] = ~16'b0;
    assign data[165] = ~16'b0;
    assign data[166] = ~16'b0;
    assign data[167] = ~16'b0;
    assign data[168] = ~16'b0;
    assign data[169] = ~16'b0;
    assign data[170] = 16'b0;
    assign data[171] = 16'b0;
    assign data[172] = ~16'b0;
    assign data[173] = ~16'b0;
    assign data[174] = ~16'b0;
    assign data[175] = ~16'b0;
    assign data[176] = ~16'b0;
    assign data[177] = ~16'b0;
    assign data[178] = ~16'b0;
    assign data[179] = ~16'b0;
    assign data[180] = 16'b0;
    assign data[181] = 16'b0;
    assign data[182] = ~16'b0;
    assign data[183] = ~16'b0;
    assign data[184] = ~16'b0;
    assign data[185] = ~16'b0;
    assign data[186] = ~16'b0;
    assign data[187] = ~16'b0;
    assign data[188] = ~16'b0;
    assign data[189] = ~16'b0;
    assign data[190] = 16'b0;
    assign data[191] = 16'b0;
    assign data[192] = ~16'b0;
    assign data[193] = ~16'b0;
    assign data[194] = ~16'b0;
    assign data[195] = ~16'b0;
    assign data[196] = ~16'b0;
    assign data[197] = ~16'b0;
    assign data[198] = ~16'b0;
    assign data[199] = ~16'b0;
    assign data[200] = 16'b0;
    assign data[201] = 16'b0;
    assign data[202] = ~16'b0;
    assign data[203] = ~16'b0;
    assign data[204] = ~16'b0;
    assign data[205] = ~16'b0;
    assign data[206] = ~16'b0;
    assign data[207] = ~16'b0;
    assign data[208] = ~16'b0;
    assign data[209] = ~16'b0;
    assign data[210] = 16'b0;
    assign data[211] = 16'b0;
    assign data[212] = ~16'b0;
    assign data[213] = ~16'b0;
    assign data[214] = ~16'b0;
    assign data[215] = ~16'b0;
    assign data[216] = ~16'b0;
    assign data[217] = ~16'b0;
    assign data[218] = ~16'b0;
    assign data[219] = ~16'b0;
    assign data[220] = 16'b0;
    assign data[221] = 16'b0;
    assign data[222] = ~16'b0;
    assign data[223] = ~16'b0;
    assign data[224] = ~16'b0;
    assign data[225] = ~16'b0;
    assign data[226] = ~16'b0;
    assign data[227] = ~16'b0;
    assign data[228] = ~16'b0;
    assign data[229] = ~16'b0;
    assign data[230] = 16'b0;
    assign data[231] = 16'b0;
    assign data[232] = ~16'b0;
    assign data[233] = ~16'b0;
    assign data[234] = ~16'b0;
    assign data[235] = ~16'b0;
    assign data[236] = ~16'b0;
    assign data[237] = ~16'b0;
    assign data[238] = ~16'b0;
    assign data[239] = ~16'b0;
    assign data[240] = 16'b0;
    assign data[241] = 16'b0;
    assign data[242] = ~16'b0;
    assign data[243] = ~16'b0;
    assign data[244] = ~16'b0;
    assign data[245] = ~16'b0;
    assign data[246] = ~16'b0;
    assign data[247] = ~16'b0;
    assign data[248] = ~16'b0;
    assign data[249] = ~16'b0;
    assign data[250] = 16'b0;
    assign data[251] = 16'b0;
    assign data[252] = ~16'b0;
    assign data[253] = ~16'b0;
    assign data[254] = ~16'b0;
    assign data[255] = ~16'b0;
    assign data[256] = ~16'b0;
    assign data[257] = ~16'b0;
    assign data[258] = ~16'b0;
    assign data[259] = ~16'b0;
    assign data[260] = 16'b0;
    assign data[261] = 16'b0;
    assign data[262] = ~16'b0;
    assign data[263] = ~16'b0;
    assign data[264] = ~16'b0;
    assign data[265] = ~16'b0;
    assign data[266] = ~16'b0;
    assign data[267] = ~16'b0;
    assign data[268] = ~16'b0;
    assign data[269] = ~16'b0;
    assign data[270] = 16'b0;
    assign data[271] = 16'b0;
    assign data[272] = ~16'b0;
    assign data[273] = ~16'b0;
    assign data[274] = ~16'b0;
    assign data[275] = ~16'b0;
    assign data[276] = ~16'b0;
    assign data[277] = ~16'b0;
    assign data[278] = ~16'b0;
    assign data[279] = ~16'b0;
    assign data[280] = 16'b0;
    assign data[281] = 16'b0;
    assign data[282] = 16'b0;
    assign data[283] = 16'b0;
    assign data[284] = 16'b0;
    assign data[285] = 16'b0;
    assign data[286] = 16'b0;
    assign data[287] = 16'b0;
    assign data[288] = 16'b0;
    assign data[289] = 16'b0;
    assign data[290] = 16'b0;
    assign data[291] = 16'b0;
    assign data[292] = 16'b0;
    assign data[293] = 16'b0;
    assign data[294] = 16'b0;
    assign data[295] = 16'b0;
    assign data[296] = 16'b0;
    assign data[297] = 16'b0;
    assign data[298] = 16'b0;
    assign data[299] = 16'b0;
    assign data[300] = ~16'b0;
    assign data[301] = ~16'b0;
    assign data[302] = ~16'b0;
    assign data[303] = ~16'b0;
    assign data[304] = ~16'b0;
    assign data[305] = ~16'b0;
    assign data[306] = ~16'b0;
    assign data[307] = ~16'b0;
    assign data[308] = ~16'b0;
    assign data[309] = ~16'b0;
    assign data[310] = ~16'b0;
    assign data[311] = ~16'b0;
    assign data[312] = ~16'b0;
    assign data[313] = ~16'b0;
    assign data[314] = ~16'b0;
    assign data[315] = ~16'b0;
    assign data[316] = ~16'b0;
    assign data[317] = ~16'b0;
    assign data[318] = ~16'b0;
    assign data[319] = ~16'b0;
    assign data[320] = ~16'b0;
    assign data[321] = ~16'b0;
    assign data[322] = ~16'b0;
    assign data[323] = ~16'b0;
    assign data[324] = ~16'b0;
    assign data[325] = ~16'b0;
    assign data[326] = ~16'b0;
    assign data[327] = ~16'b0;
    assign data[328] = ~16'b0;
    assign data[329] = ~16'b0;
    assign data[330] = ~16'b0;
    assign data[331] = ~16'b0;
    assign data[332] = ~16'b0;
    assign data[333] = ~16'b0;
    assign data[334] = ~16'b0;
    assign data[335] = ~16'b0;
    assign data[336] = ~16'b0;
    assign data[337] = ~16'b0;
    assign data[338] = ~16'b0;
    assign data[339] = ~16'b0;
    assign data[340] = ~16'b0;
    assign data[341] = ~16'b0;
    assign data[342] = ~16'b0;
    assign data[343] = ~16'b0;
    assign data[344] = ~16'b0;
    assign data[345] = ~16'b0;
    assign data[346] = ~16'b0;
    assign data[347] = ~16'b0;
    assign data[348] = ~16'b0;
    assign data[349] = ~16'b0;
    assign data[350] = ~16'b0;
    assign data[351] = ~16'b0;
    assign data[352] = ~16'b0;
    assign data[353] = ~16'b0;
    assign data[354] = ~16'b0;
    assign data[355] = ~16'b0;
    assign data[356] = ~16'b0;
    assign data[357] = ~16'b0;
    assign data[358] = ~16'b0;
    assign data[359] = ~16'b0;
    assign data[360] = ~16'b0;
    assign data[361] = ~16'b0;
    assign data[362] = ~16'b0;
    assign data[363] = ~16'b0;
    assign data[364] = ~16'b0;
    assign data[365] = ~16'b0;
    assign data[366] = ~16'b0;
    assign data[367] = ~16'b0;
    assign data[368] = ~16'b0;
    assign data[369] = ~16'b0;
    assign data[370] = ~16'b0;
    assign data[371] = ~16'b0;
    assign data[372] = ~16'b0;
    assign data[373] = ~16'b0;
    assign data[374] = ~16'b0;
    assign data[375] = ~16'b0;
    assign data[376] = ~16'b0;
    assign data[377] = ~16'b0;
    assign data[378] = ~16'b0;
    assign data[379] = ~16'b0;
    assign data[380] = ~16'b0;
    assign data[381] = ~16'b0;
    assign data[382] = ~16'b0;
    assign data[383] = ~16'b0;
    assign data[384] = ~16'b0;
    assign data[385] = ~16'b0;
    assign data[386] = ~16'b0;
    assign data[387] = ~16'b0;
    assign data[388] = ~16'b0;
    assign data[389] = ~16'b0;
    assign data[390] = ~16'b0;
    assign data[391] = ~16'b0;
    assign data[392] = ~16'b0;
    assign data[393] = ~16'b0;
    assign data[394] = ~16'b0;
    assign data[395] = ~16'b0;
    assign data[396] = ~16'b0;
    assign data[397] = ~16'b0;
    assign data[398] = ~16'b0;
    assign data[399] = ~16'b0;
    assign data[400] = 16'b0;
    assign data[401] = 16'b0;
    assign data[402] = 16'b0;
    assign data[403] = 16'b0;
    assign data[404] = 16'b0;
    assign data[405] = 16'b0;
    assign data[406] = 16'b0;
    assign data[407] = 16'b0;
    assign data[408] = 16'b0;
    assign data[409] = 16'b0;
    assign data[410] = 16'b0;
    assign data[411] = 16'b0;
    assign data[412] = 16'b0;
    assign data[413] = 16'b0;
    assign data[414] = 16'b0;
    assign data[415] = 16'b0;
    assign data[416] = 16'b0;
    assign data[417] = 16'b0;
    assign data[418] = 16'b0;
    assign data[419] = 16'b0;
    assign data[420] = 16'b0;
    assign data[421] = 16'b0;
    assign data[422] = ~16'b0;
    assign data[423] = ~16'b0;
    assign data[424] = ~16'b0;
    assign data[425] = ~16'b0;
    assign data[426] = ~16'b0;
    assign data[427] = ~16'b0;
    assign data[428] = ~16'b0;
    assign data[429] = ~16'b0;
    assign data[430] = 16'b0;
    assign data[431] = 16'b0;
    assign data[432] = ~16'b0;
    assign data[433] = ~16'b0;
    assign data[434] = ~16'b0;
    assign data[435] = ~16'b0;
    assign data[436] = ~16'b0;
    assign data[437] = ~16'b0;
    assign data[438] = ~16'b0;
    assign data[439] = ~16'b0;
    assign data[440] = 16'b0;
    assign data[441] = 16'b0;
    assign data[442] = ~16'b0;
    assign data[443] = ~16'b0;
    assign data[444] = ~16'b0;
    assign data[445] = ~16'b0;
    assign data[446] = ~16'b0;
    assign data[447] = ~16'b0;
    assign data[448] = ~16'b0;
    assign data[449] = ~16'b0;
    assign data[450] = 16'b0;
    assign data[451] = 16'b0;
    assign data[452] = ~16'b0;
    assign data[453] = ~16'b0;
    assign data[454] = ~16'b0;
    assign data[455] = ~16'b0;
    assign data[456] = ~16'b0;
    assign data[457] = ~16'b0;
    assign data[458] = ~16'b0;
    assign data[459] = ~16'b0;
    assign data[460] = 16'b0;
    assign data[461] = 16'b0;
    assign data[462] = ~16'b0;
    assign data[463] = ~16'b0;
    assign data[464] = ~16'b0;
    assign data[465] = ~16'b0;
    assign data[466] = ~16'b0;
    assign data[467] = ~16'b0;
    assign data[468] = ~16'b0;
    assign data[469] = ~16'b0;
    assign data[470] = 16'b0;
    assign data[471] = 16'b0;
    assign data[472] = ~16'b0;
    assign data[473] = ~16'b0;
    assign data[474] = ~16'b0;
    assign data[475] = ~16'b0;
    assign data[476] = ~16'b0;
    assign data[477] = ~16'b0;
    assign data[478] = ~16'b0;
    assign data[479] = ~16'b0;
    assign data[480] = 16'b0;
    assign data[481] = 16'b0;
    assign data[482] = ~16'b0;
    assign data[483] = ~16'b0;
    assign data[484] = ~16'b0;
    assign data[485] = ~16'b0;
    assign data[486] = ~16'b0;
    assign data[487] = ~16'b0;
    assign data[488] = ~16'b0;
    assign data[489] = ~16'b0;
    assign data[490] = 16'b0;
    assign data[491] = 16'b0;
    assign data[492] = ~16'b0;
    assign data[493] = ~16'b0;
    assign data[494] = ~16'b0;
    assign data[495] = ~16'b0;
    assign data[496] = ~16'b0;
    assign data[497] = ~16'b0;
    assign data[498] = ~16'b0;
    assign data[499] = ~16'b0;
    assign data[500] = 16'b0;
    assign data[501] = 16'b0;
    assign data[502] = ~16'b0;
    assign data[503] = ~16'b0;
    assign data[504] = ~16'b0;
    assign data[505] = ~16'b0;
    assign data[506] = ~16'b0;
    assign data[507] = ~16'b0;
    assign data[508] = ~16'b0;
    assign data[509] = ~16'b0;
    assign data[510] = 16'b0;
    assign data[511] = 16'b0;
    assign data[512] = ~16'b0;
    assign data[513] = ~16'b0;
    assign data[514] = ~16'b0;
    assign data[515] = ~16'b0;
    assign data[516] = ~16'b0;
    assign data[517] = ~16'b0;
    assign data[518] = ~16'b0;
    assign data[519] = ~16'b0;
    assign data[520] = 16'b0;
    assign data[521] = 16'b0;
    assign data[522] = ~16'b0;
    assign data[523] = ~16'b0;
    assign data[524] = ~16'b0;
    assign data[525] = ~16'b0;
    assign data[526] = ~16'b0;
    assign data[527] = ~16'b0;
    assign data[528] = ~16'b0;
    assign data[529] = ~16'b0;
    assign data[530] = 16'b0;
    assign data[531] = 16'b0;
    assign data[532] = ~16'b0;
    assign data[533] = ~16'b0;
    assign data[534] = ~16'b0;
    assign data[535] = ~16'b0;
    assign data[536] = ~16'b0;
    assign data[537] = ~16'b0;
    assign data[538] = ~16'b0;
    assign data[539] = ~16'b0;
    assign data[540] = 16'b0;
    assign data[541] = 16'b0;
    assign data[542] = ~16'b0;
    assign data[543] = ~16'b0;
    assign data[544] = ~16'b0;
    assign data[545] = ~16'b0;
    assign data[546] = ~16'b0;
    assign data[547] = ~16'b0;
    assign data[548] = ~16'b0;
    assign data[549] = ~16'b0;
    assign data[550] = 16'b0;
    assign data[551] = 16'b0;
    assign data[552] = ~16'b0;
    assign data[553] = ~16'b0;
    assign data[554] = ~16'b0;
    assign data[555] = ~16'b0;
    assign data[556] = ~16'b0;
    assign data[557] = ~16'b0;
    assign data[558] = ~16'b0;
    assign data[559] = ~16'b0;
    assign data[560] = 16'b0;
    assign data[561] = 16'b0;
    assign data[562] = ~16'b0;
    assign data[563] = ~16'b0;
    assign data[564] = ~16'b0;
    assign data[565] = ~16'b0;
    assign data[566] = ~16'b0;
    assign data[567] = ~16'b0;
    assign data[568] = ~16'b0;
    assign data[569] = ~16'b0;
    assign data[570] = 16'b0;
    assign data[571] = 16'b0;
    assign data[572] = ~16'b0;
    assign data[573] = ~16'b0;
    assign data[574] = ~16'b0;
    assign data[575] = ~16'b0;
    assign data[576] = ~16'b0;
    assign data[577] = ~16'b0;
    assign data[578] = ~16'b0;
    assign data[579] = ~16'b0;
    assign data[580] = 16'b0;
    assign data[581] = 16'b0;
    assign data[582] = ~16'b0;
    assign data[583] = ~16'b0;
    assign data[584] = ~16'b0;
    assign data[585] = ~16'b0;
    assign data[586] = ~16'b0;
    assign data[587] = ~16'b0;
    assign data[588] = ~16'b0;
    assign data[589] = ~16'b0;
    assign data[590] = 16'b0;
    assign data[591] = 16'b0;
    assign data[592] = ~16'b0;
    assign data[593] = ~16'b0;
    assign data[594] = ~16'b0;
    assign data[595] = ~16'b0;
    assign data[596] = ~16'b0;
    assign data[597] = ~16'b0;
    assign data[598] = ~16'b0;
    assign data[599] = ~16'b0;
    assign data[600] = 16'b0;
    assign data[601] = 16'b0;
    assign data[602] = ~16'b0;
    assign data[603] = ~16'b0;
    assign data[604] = ~16'b0;
    assign data[605] = ~16'b0;
    assign data[606] = ~16'b0;
    assign data[607] = ~16'b0;
    assign data[608] = ~16'b0;
    assign data[609] = ~16'b0;
    assign data[610] = 16'b0;
    assign data[611] = 16'b0;
    assign data[612] = ~16'b0;
    assign data[613] = ~16'b0;
    assign data[614] = ~16'b0;
    assign data[615] = ~16'b0;
    assign data[616] = ~16'b0;
    assign data[617] = ~16'b0;
    assign data[618] = ~16'b0;
    assign data[619] = ~16'b0;
    assign data[620] = 16'b0;
    assign data[621] = 16'b0;
    assign data[622] = ~16'b0;
    assign data[623] = ~16'b0;
    assign data[624] = ~16'b0;
    assign data[625] = ~16'b0;
    assign data[626] = ~16'b0;
    assign data[627] = ~16'b0;
    assign data[628] = ~16'b0;
    assign data[629] = ~16'b0;
    assign data[630] = 16'b0;
    assign data[631] = 16'b0;
    assign data[632] = ~16'b0;
    assign data[633] = ~16'b0;
    assign data[634] = ~16'b0;
    assign data[635] = ~16'b0;
    assign data[636] = ~16'b0;
    assign data[637] = ~16'b0;
    assign data[638] = ~16'b0;
    assign data[639] = ~16'b0;
    assign data[640] = 16'b0;
    assign data[641] = 16'b0;
    assign data[642] = ~16'b0;
    assign data[643] = ~16'b0;
    assign data[644] = ~16'b0;
    assign data[645] = ~16'b0;
    assign data[646] = ~16'b0;
    assign data[647] = ~16'b0;
    assign data[648] = ~16'b0;
    assign data[649] = ~16'b0;
    assign data[650] = 16'b0;
    assign data[651] = 16'b0;
    assign data[652] = ~16'b0;
    assign data[653] = ~16'b0;
    assign data[654] = ~16'b0;
    assign data[655] = ~16'b0;
    assign data[656] = ~16'b0;
    assign data[657] = ~16'b0;
    assign data[658] = ~16'b0;
    assign data[659] = ~16'b0;
    assign data[660] = 16'b0;
    assign data[661] = 16'b0;
    assign data[662] = ~16'b0;
    assign data[663] = ~16'b0;
    assign data[664] = ~16'b0;
    assign data[665] = ~16'b0;
    assign data[666] = ~16'b0;
    assign data[667] = ~16'b0;
    assign data[668] = ~16'b0;
    assign data[669] = ~16'b0;
    assign data[670] = 16'b0;
    assign data[671] = 16'b0;
    assign data[672] = ~16'b0;
    assign data[673] = ~16'b0;
    assign data[674] = ~16'b0;
    assign data[675] = ~16'b0;
    assign data[676] = ~16'b0;
    assign data[677] = ~16'b0;
    assign data[678] = ~16'b0;
    assign data[679] = ~16'b0;
    assign data[680] = 16'b0;
    assign data[681] = 16'b0;
    assign data[682] = ~16'b0;
    assign data[683] = ~16'b0;
    assign data[684] = ~16'b0;
    assign data[685] = ~16'b0;
    assign data[686] = ~16'b0;
    assign data[687] = ~16'b0;
    assign data[688] = ~16'b0;
    assign data[689] = ~16'b0;
    assign data[690] = 16'b0;
    assign data[691] = 16'b0;
    assign data[692] = ~16'b0;
    assign data[693] = ~16'b0;
    assign data[694] = ~16'b0;
    assign data[695] = ~16'b0;
    assign data[696] = ~16'b0;
    assign data[697] = ~16'b0;
    assign data[698] = ~16'b0;
    assign data[699] = ~16'b0;
    assign data[700] = 16'b0;
    assign data[701] = 16'b0;
    assign data[702] = ~16'b0;
    assign data[703] = ~16'b0;
    assign data[704] = ~16'b0;
    assign data[705] = ~16'b0;
    assign data[706] = ~16'b0;
    assign data[707] = ~16'b0;
    assign data[708] = ~16'b0;
    assign data[709] = ~16'b0;
    assign data[710] = 16'b0;
    assign data[711] = 16'b0;
    assign data[712] = 16'b0;
    assign data[713] = 16'b0;
    assign data[714] = 16'b0;
    assign data[715] = 16'b0;
    assign data[716] = 16'b0;
    assign data[717] = 16'b0;
    assign data[718] = 16'b0;
    assign data[719] = 16'b0;
    assign data[720] = 16'b0;
    assign data[721] = 16'b0;
    assign data[722] = 16'b0;
    assign data[723] = 16'b0;
    assign data[724] = 16'b0;
    assign data[725] = 16'b0;
    assign data[726] = 16'b0;
    assign data[727] = 16'b0;
    assign data[728] = 16'b0;
    assign data[729] = 16'b0;
    assign data[730] = ~16'b0;
    assign data[731] = ~16'b0;
    assign data[732] = ~16'b0;
    assign data[733] = ~16'b0;
    assign data[734] = ~16'b0;
    assign data[735] = ~16'b0;
    assign data[736] = ~16'b0;
    assign data[737] = ~16'b0;
    assign data[738] = ~16'b0;
    assign data[739] = ~16'b0;
    assign data[740] = ~16'b0;
    assign data[741] = ~16'b0;
    assign data[742] = ~16'b0;
    assign data[743] = ~16'b0;
    assign data[744] = ~16'b0;
    assign data[745] = ~16'b0;
    assign data[746] = ~16'b0;
    assign data[747] = ~16'b0;
    assign data[748] = ~16'b0;
    assign data[749] = ~16'b0;
    assign data[750] = ~16'b0;
    assign data[751] = ~16'b0;
    assign data[752] = ~16'b0;
    assign data[753] = ~16'b0;
    assign data[754] = ~16'b0;
    assign data[755] = ~16'b0;
    assign data[756] = ~16'b0;
    assign data[757] = ~16'b0;
    assign data[758] = ~16'b0;
    assign data[759] = ~16'b0;
    assign data[760] = ~16'b0;
    assign data[761] = ~16'b0;
    assign data[762] = ~16'b0;
    assign data[763] = ~16'b0;
    assign data[764] = ~16'b0;
    assign data[765] = ~16'b0;
    assign data[766] = ~16'b0;
    assign data[767] = ~16'b0;
    assign data[768] = ~16'b0;
    assign data[769] = ~16'b0;
    assign data[770] = ~16'b0;
    assign data[771] = ~16'b0;
    assign data[772] = ~16'b0;
    assign data[773] = ~16'b0;
    assign data[774] = ~16'b0;
    assign data[775] = ~16'b0;
    assign data[776] = ~16'b0;
    assign data[777] = ~16'b0;
    assign data[778] = ~16'b0;
    assign data[779] = ~16'b0;
    assign data[780] = ~16'b0;
    assign data[781] = ~16'b0;
    assign data[782] = ~16'b0;
    assign data[783] = ~16'b0;
    assign data[784] = ~16'b0;
    assign data[785] = ~16'b0;
    assign data[786] = ~16'b0;
    assign data[787] = ~16'b0;
    assign data[788] = ~16'b0;
    assign data[789] = ~16'b0;
    assign data[790] = ~16'b0;
    assign data[791] = ~16'b0;
    assign data[792] = ~16'b0;
    assign data[793] = ~16'b0;
    assign data[794] = ~16'b0;
    assign data[795] = ~16'b0;
    assign data[796] = ~16'b0;
    assign data[797] = ~16'b0;
    assign data[798] = ~16'b0;
    assign data[799] = ~16'b0;
    assign data[800] = ~16'b0;
    assign data[801] = ~16'b0;
    assign data[802] = ~16'b0;
    assign data[803] = ~16'b0;
    assign data[804] = ~16'b0;
    assign data[805] = ~16'b0;
    assign data[806] = ~16'b0;
    assign data[807] = ~16'b0;
    assign data[808] = ~16'b0;
    assign data[809] = ~16'b0;
    assign data[810] = ~16'b0;
    assign data[811] = ~16'b0;
    assign data[812] = ~16'b0;
    assign data[813] = ~16'b0;
    assign data[814] = ~16'b0;
    assign data[815] = ~16'b0;
    assign data[816] = ~16'b0;
    assign data[817] = ~16'b0;
    assign data[818] = ~16'b0;
    assign data[819] = ~16'b0;
    assign data[820] = ~16'b0;
    assign data[821] = ~16'b0;
    assign data[822] = ~16'b0;
    assign data[823] = ~16'b0;
    assign data[824] = ~16'b0;
    assign data[825] = ~16'b0;
    assign data[826] = ~16'b0;
    assign data[827] = ~16'b0;
    assign data[828] = ~16'b0;
    assign data[829] = ~16'b0;
    assign data[830] = ~16'b0;
    assign data[831] = ~16'b0;
    assign data[832] = ~16'b0;
    assign data[833] = ~16'b0;
    assign data[834] = ~16'b0;
    assign data[835] = ~16'b0;
    assign data[836] = ~16'b0;
    assign data[837] = ~16'b0;
    assign data[838] = ~16'b0;
    assign data[839] = ~16'b0;
    assign data[840] = ~16'b0;
    assign data[841] = ~16'b0;
    assign data[842] = ~16'b0;
    assign data[843] = ~16'b0;
    assign data[844] = ~16'b0;
    assign data[845] = ~16'b0;
    assign data[846] = ~16'b0;
    assign data[847] = ~16'b0;
    assign data[848] = ~16'b0;
    assign data[849] = ~16'b0;
    assign data[850] = ~16'b0;
    assign data[851] = ~16'b0;
    assign data[852] = ~16'b0;
    assign data[853] = ~16'b0;
    assign data[854] = ~16'b0;
    assign data[855] = ~16'b0;
    assign data[856] = ~16'b0;
    assign data[857] = ~16'b0;
    assign data[858] = ~16'b0;
    assign data[859] = ~16'b0;
    assign data[860] = ~16'b0;
    assign data[861] = ~16'b0;
    assign data[862] = ~16'b0;
    assign data[863] = ~16'b0;
    assign data[864] = ~16'b0;
    assign data[865] = ~16'b0;
    assign data[866] = ~16'b0;
    assign data[867] = ~16'b0;
    assign data[868] = ~16'b0;
    assign data[869] = ~16'b0;
    assign data[870] = ~16'b0;
    assign data[871] = ~16'b0;
    assign data[872] = ~16'b0;
    assign data[873] = ~16'b0;
    assign data[874] = ~16'b0;
    assign data[875] = ~16'b0;
    assign data[876] = ~16'b0;
    assign data[877] = ~16'b0;
    assign data[878] = ~16'b0;
    assign data[879] = ~16'b0;
    assign data[880] = ~16'b0;
    assign data[881] = ~16'b0;
    assign data[882] = ~16'b0;
    assign data[883] = ~16'b0;
    assign data[884] = ~16'b0;
    assign data[885] = ~16'b0;
    assign data[886] = ~16'b0;
    assign data[887] = ~16'b0;
    assign data[888] = ~16'b0;
    assign data[889] = ~16'b0;
    assign data[890] = ~16'b0;
    assign data[891] = ~16'b0;
    assign data[892] = ~16'b0;
    assign data[893] = ~16'b0;
    assign data[894] = ~16'b0;
    assign data[895] = ~16'b0;
    assign data[896] = ~16'b0;
    assign data[897] = ~16'b0;
    assign data[898] = ~16'b0;
    assign data[899] = ~16'b0;
    assign data[900] = ~16'b0;
    assign data[901] = ~16'b0;
    assign data[902] = ~16'b0;
    assign data[903] = ~16'b0;
    assign data[904] = ~16'b0;
    assign data[905] = ~16'b0;
    assign data[906] = ~16'b0;
    assign data[907] = ~16'b0;
    assign data[908] = ~16'b0;
    assign data[909] = ~16'b0;
    assign data[910] = ~16'b0;
    assign data[911] = ~16'b0;
    assign data[912] = ~16'b0;
    assign data[913] = ~16'b0;
    assign data[914] = ~16'b0;
    assign data[915] = ~16'b0;
    assign data[916] = ~16'b0;
    assign data[917] = ~16'b0;
    assign data[918] = ~16'b0;
    assign data[919] = ~16'b0;
    assign data[920] = ~16'b0;
    assign data[921] = ~16'b0;
    assign data[922] = ~16'b0;
    assign data[923] = ~16'b0;
    assign data[924] = ~16'b0;
    assign data[925] = ~16'b0;
    assign data[926] = ~16'b0;
    assign data[927] = ~16'b0;
    assign data[928] = ~16'b0;
    assign data[929] = ~16'b0;
    assign data[930] = 16'b0;
    assign data[931] = 16'b0;
    assign data[932] = 16'b0;
    assign data[933] = 16'b0;
    assign data[934] = 16'b0;
    assign data[935] = 16'b0;
    assign data[936] = 16'b0;
    assign data[937] = 16'b0;
    assign data[938] = 16'b0;
    assign data[939] = 16'b0;
    assign data[940] = 16'b0;
    assign data[941] = 16'b0;
    assign data[942] = 16'b0;
    assign data[943] = 16'b0;
    assign data[944] = 16'b0;
    assign data[945] = 16'b0;
    assign data[946] = 16'b0;
    assign data[947] = 16'b0;
    assign data[948] = 16'b0;
    assign data[949] = 16'b0;
    assign data[950] = 16'b0;
    assign data[951] = 16'b0;
    assign data[952] = ~16'b0;
    assign data[953] = ~16'b0;
    assign data[954] = ~16'b0;
    assign data[955] = ~16'b0;
    assign data[956] = ~16'b0;
    assign data[957] = ~16'b0;
    assign data[958] = ~16'b0;
    assign data[959] = ~16'b0;
    assign data[960] = 16'b0;
    assign data[961] = 16'b0;
    assign data[962] = ~16'b0;
    assign data[963] = ~16'b0;
    assign data[964] = ~16'b0;
    assign data[965] = ~16'b0;
    assign data[966] = ~16'b0;
    assign data[967] = ~16'b0;
    assign data[968] = ~16'b0;
    assign data[969] = ~16'b0;
    assign data[970] = 16'b0;
    assign data[971] = 16'b0;
    assign data[972] = ~16'b0;
    assign data[973] = ~16'b0;
    assign data[974] = ~16'b0;
    assign data[975] = ~16'b0;
    assign data[976] = ~16'b0;
    assign data[977] = ~16'b0;
    assign data[978] = ~16'b0;
    assign data[979] = ~16'b0;
    assign data[980] = 16'b0;
    assign data[981] = 16'b0;
    assign data[982] = ~16'b0;
    assign data[983] = ~16'b0;
    assign data[984] = ~16'b0;
    assign data[985] = ~16'b0;
    assign data[986] = ~16'b0;
    assign data[987] = ~16'b0;
    assign data[988] = ~16'b0;
    assign data[989] = ~16'b0;
    assign data[990] = 16'b0;
    assign data[991] = 16'b0;
    assign data[992] = ~16'b0;
    assign data[993] = ~16'b0;
    assign data[994] = ~16'b0;
    assign data[995] = ~16'b0;
    assign data[996] = ~16'b0;
    assign data[997] = ~16'b0;
    assign data[998] = ~16'b0;
    assign data[999] = ~16'b0;
    assign data[1000] = 16'b0;
    assign data[1001] = 16'b0;
    assign data[1002] = ~16'b0;
    assign data[1003] = ~16'b0;
    assign data[1004] = ~16'b0;
    assign data[1005] = ~16'b0;
    assign data[1006] = ~16'b0;
    assign data[1007] = ~16'b0;
    assign data[1008] = ~16'b0;
    assign data[1009] = ~16'b0;
    assign data[1010] = 16'b0;
    assign data[1011] = 16'b0;
    assign data[1012] = ~16'b0;
    assign data[1013] = ~16'b0;
    assign data[1014] = ~16'b0;
    assign data[1015] = ~16'b0;
    assign data[1016] = ~16'b0;
    assign data[1017] = ~16'b0;
    assign data[1018] = ~16'b0;
    assign data[1019] = ~16'b0;
    assign data[1020] = 16'b0;
    assign data[1021] = 16'b0;
    assign data[1022] = ~16'b0;
    assign data[1023] = ~16'b0;
    assign data[1024] = ~16'b0;
    assign data[1025] = ~16'b0;
    assign data[1026] = ~16'b0;
    assign data[1027] = ~16'b0;
    assign data[1028] = ~16'b0;
    assign data[1029] = ~16'b0;
    assign data[1030] = 16'b0;
    assign data[1031] = 16'b0;
    assign data[1032] = ~16'b0;
    assign data[1033] = ~16'b0;
    assign data[1034] = ~16'b0;
    assign data[1035] = ~16'b0;
    assign data[1036] = ~16'b0;
    assign data[1037] = ~16'b0;
    assign data[1038] = ~16'b0;
    assign data[1039] = ~16'b0;
    assign data[1040] = 16'b0;
    assign data[1041] = 16'b0;
    assign data[1042] = ~16'b0;
    assign data[1043] = ~16'b0;
    assign data[1044] = ~16'b0;
    assign data[1045] = ~16'b0;
    assign data[1046] = ~16'b0;
    assign data[1047] = ~16'b0;
    assign data[1048] = ~16'b0;
    assign data[1049] = ~16'b0;
    assign data[1050] = 16'b0;
    assign data[1051] = 16'b0;
    assign data[1052] = ~16'b0;
    assign data[1053] = ~16'b0;
    assign data[1054] = ~16'b0;
    assign data[1055] = ~16'b0;
    assign data[1056] = ~16'b0;
    assign data[1057] = ~16'b0;
    assign data[1058] = ~16'b0;
    assign data[1059] = ~16'b0;
    assign data[1060] = 16'b0;
    assign data[1061] = 16'b0;
    assign data[1062] = ~16'b0;
    assign data[1063] = ~16'b0;
    assign data[1064] = ~16'b0;
    assign data[1065] = ~16'b0;
    assign data[1066] = ~16'b0;
    assign data[1067] = ~16'b0;
    assign data[1068] = ~16'b0;
    assign data[1069] = ~16'b0;
    assign data[1070] = 16'b0;
    assign data[1071] = 16'b0;
    assign data[1072] = ~16'b0;
    assign data[1073] = ~16'b0;
    assign data[1074] = ~16'b0;
    assign data[1075] = ~16'b0;
    assign data[1076] = ~16'b0;
    assign data[1077] = ~16'b0;
    assign data[1078] = ~16'b0;
    assign data[1079] = ~16'b0;
    assign data[1080] = 16'b0;
    assign data[1081] = 16'b0;
    assign data[1082] = ~16'b0;
    assign data[1083] = ~16'b0;
    assign data[1084] = ~16'b0;
    assign data[1085] = ~16'b0;
    assign data[1086] = ~16'b0;
    assign data[1087] = ~16'b0;
    assign data[1088] = ~16'b0;
    assign data[1089] = ~16'b0;
    assign data[1090] = 16'b0;
    assign data[1091] = 16'b0;
    assign data[1092] = ~16'b0;
    assign data[1093] = ~16'b0;
    assign data[1094] = ~16'b0;
    assign data[1095] = ~16'b0;
    assign data[1096] = ~16'b0;
    assign data[1097] = ~16'b0;
    assign data[1098] = ~16'b0;
    assign data[1099] = ~16'b0;
    assign data[1100] = 16'b0;
    assign data[1101] = 16'b0;
    assign data[1102] = ~16'b0;
    assign data[1103] = ~16'b0;
    assign data[1104] = ~16'b0;
    assign data[1105] = ~16'b0;
    assign data[1106] = ~16'b0;
    assign data[1107] = ~16'b0;
    assign data[1108] = ~16'b0;
    assign data[1109] = ~16'b0;
    assign data[1110] = 16'b0;
    assign data[1111] = 16'b0;
    assign data[1112] = ~16'b0;
    assign data[1113] = ~16'b0;
    assign data[1114] = ~16'b0;
    assign data[1115] = ~16'b0;
    assign data[1116] = ~16'b0;
    assign data[1117] = ~16'b0;
    assign data[1118] = ~16'b0;
    assign data[1119] = ~16'b0;
    assign data[1120] = 16'b0;
    assign data[1121] = 16'b0;
    assign data[1122] = ~16'b0;
    assign data[1123] = ~16'b0;
    assign data[1124] = ~16'b0;
    assign data[1125] = ~16'b0;
    assign data[1126] = ~16'b0;
    assign data[1127] = ~16'b0;
    assign data[1128] = ~16'b0;
    assign data[1129] = ~16'b0;
    assign data[1130] = 16'b0;
    assign data[1131] = 16'b0;
    assign data[1132] = ~16'b0;
    assign data[1133] = ~16'b0;
    assign data[1134] = ~16'b0;
    assign data[1135] = ~16'b0;
    assign data[1136] = ~16'b0;
    assign data[1137] = ~16'b0;
    assign data[1138] = ~16'b0;
    assign data[1139] = ~16'b0;
    assign data[1140] = 16'b0;
    assign data[1141] = 16'b0;
    assign data[1142] = ~16'b0;
    assign data[1143] = ~16'b0;
    assign data[1144] = ~16'b0;
    assign data[1145] = ~16'b0;
    assign data[1146] = ~16'b0;
    assign data[1147] = ~16'b0;
    assign data[1148] = ~16'b0;
    assign data[1149] = ~16'b0;
    assign data[1150] = 16'b0;
    assign data[1151] = 16'b0;
    assign data[1152] = ~16'b0;
    assign data[1153] = ~16'b0;
    assign data[1154] = ~16'b0;
    assign data[1155] = ~16'b0;
    assign data[1156] = ~16'b0;
    assign data[1157] = ~16'b0;
    assign data[1158] = ~16'b0;
    assign data[1159] = ~16'b0;
    assign data[1160] = 16'b0;
    assign data[1161] = 16'b0;
    assign data[1162] = ~16'b0;
    assign data[1163] = ~16'b0;
    assign data[1164] = ~16'b0;
    assign data[1165] = ~16'b0;
    assign data[1166] = ~16'b0;
    assign data[1167] = ~16'b0;
    assign data[1168] = ~16'b0;
    assign data[1169] = ~16'b0;
    assign data[1170] = 16'b0;
    assign data[1171] = 16'b0;
    assign data[1172] = ~16'b0;
    assign data[1173] = ~16'b0;
    assign data[1174] = ~16'b0;
    assign data[1175] = ~16'b0;
    assign data[1176] = ~16'b0;
    assign data[1177] = ~16'b0;
    assign data[1178] = ~16'b0;
    assign data[1179] = ~16'b0;
    assign data[1180] = 16'b0;
    assign data[1181] = 16'b0;
    assign data[1182] = ~16'b0;
    assign data[1183] = ~16'b0;
    assign data[1184] = ~16'b0;
    assign data[1185] = ~16'b0;
    assign data[1186] = ~16'b0;
    assign data[1187] = ~16'b0;
    assign data[1188] = ~16'b0;
    assign data[1189] = ~16'b0;
    assign data[1190] = 16'b0;
    assign data[1191] = 16'b0;
    assign data[1192] = ~16'b0;
    assign data[1193] = ~16'b0;
    assign data[1194] = ~16'b0;
    assign data[1195] = ~16'b0;
    assign data[1196] = ~16'b0;
    assign data[1197] = ~16'b0;
    assign data[1198] = ~16'b0;
    assign data[1199] = ~16'b0;
    assign data[1200] = 16'b0;
    assign data[1201] = 16'b0;
    assign data[1202] = 16'b0;
    assign data[1203] = 16'b0;
    assign data[1204] = 16'b0;
    assign data[1205] = 16'b0;
    assign data[1206] = 16'b0;
    assign data[1207] = 16'b0;
    assign data[1208] = 16'b0;
    assign data[1209] = 16'b0;
    assign data[1210] = 16'b0;
    assign data[1211] = 16'b0;
    assign data[1212] = 16'b0;
    assign data[1213] = 16'b0;
    assign data[1214] = 16'b0;
    assign data[1215] = 16'b0;
    assign data[1216] = 16'b0;
    assign data[1217] = 16'b0;
    assign data[1218] = 16'b0;
    assign data[1219] = 16'b0;
    assign data[1220] = ~16'b0;
    assign data[1221] = ~16'b0;
    assign data[1222] = ~16'b0;
    assign data[1223] = ~16'b0;
    assign data[1224] = ~16'b0;
    assign data[1225] = ~16'b0;
    assign data[1226] = ~16'b0;
    assign data[1227] = ~16'b0;
    assign data[1228] = ~16'b0;
    assign data[1229] = ~16'b0;
    assign data[1230] = ~16'b0;
    assign data[1231] = ~16'b0;
    assign data[1232] = ~16'b0;
    assign data[1233] = ~16'b0;
    assign data[1234] = ~16'b0;
    assign data[1235] = ~16'b0;
    assign data[1236] = ~16'b0;
    assign data[1237] = ~16'b0;
    assign data[1238] = ~16'b0;
    assign data[1239] = ~16'b0;
    assign data[1240] = ~16'b0;
    assign data[1241] = ~16'b0;
    assign data[1242] = ~16'b0;
    assign data[1243] = ~16'b0;
    assign data[1244] = ~16'b0;
    assign data[1245] = ~16'b0;
    assign data[1246] = ~16'b0;
    assign data[1247] = ~16'b0;
    assign data[1248] = ~16'b0;
    assign data[1249] = ~16'b0;
    assign data[1250] = ~16'b0;
    assign data[1251] = ~16'b0;
    assign data[1252] = ~16'b0;
    assign data[1253] = ~16'b0;
    assign data[1254] = ~16'b0;
    assign data[1255] = ~16'b0;
    assign data[1256] = ~16'b0;
    assign data[1257] = ~16'b0;
    assign data[1258] = ~16'b0;
    assign data[1259] = ~16'b0;
    assign data[1260] = ~16'b0;
    assign data[1261] = ~16'b0;
    assign data[1262] = ~16'b0;
    assign data[1263] = ~16'b0;
    assign data[1264] = ~16'b0;
    assign data[1265] = ~16'b0;
    assign data[1266] = ~16'b0;
    assign data[1267] = ~16'b0;
    assign data[1268] = ~16'b0;
    assign data[1269] = ~16'b0;
    assign data[1270] = ~16'b0;
    assign data[1271] = ~16'b0;
    assign data[1272] = ~16'b0;
    assign data[1273] = ~16'b0;
    assign data[1274] = ~16'b0;
    assign data[1275] = ~16'b0;
    assign data[1276] = ~16'b0;
    assign data[1277] = ~16'b0;
    assign data[1278] = ~16'b0;
    assign data[1279] = ~16'b0;
    assign data[1280] = ~16'b0;
    assign data[1281] = ~16'b0;
    assign data[1282] = ~16'b0;
    assign data[1283] = ~16'b0;
    assign data[1284] = ~16'b0;
    assign data[1285] = ~16'b0;
    assign data[1286] = ~16'b0;
    assign data[1287] = ~16'b0;
    assign data[1288] = ~16'b0;
    assign data[1289] = ~16'b0;
    assign data[1290] = ~16'b0;
    assign data[1291] = ~16'b0;
    assign data[1292] = ~16'b0;
    assign data[1293] = ~16'b0;
    assign data[1294] = ~16'b0;
    assign data[1295] = ~16'b0;
    assign data[1296] = ~16'b0;
    assign data[1297] = ~16'b0;
    assign data[1298] = ~16'b0;
    assign data[1299] = ~16'b0;
    assign data[1300] = ~16'b0;
    assign data[1301] = ~16'b0;
    assign data[1302] = ~16'b0;
    assign data[1303] = ~16'b0;
    assign data[1304] = ~16'b0;
    assign data[1305] = ~16'b0;
    assign data[1306] = ~16'b0;
    assign data[1307] = ~16'b0;
    assign data[1308] = ~16'b0;
    assign data[1309] = ~16'b0;
    assign data[1310] = ~16'b0;
    assign data[1311] = ~16'b0;
    assign data[1312] = ~16'b0;
    assign data[1313] = ~16'b0;
    assign data[1314] = ~16'b0;
    assign data[1315] = ~16'b0;
    assign data[1316] = ~16'b0;
    assign data[1317] = ~16'b0;
    assign data[1318] = ~16'b0;
    assign data[1319] = ~16'b0;
    assign data[1320] = ~16'b0;
    assign data[1321] = ~16'b0;
    assign data[1322] = ~16'b0;
    assign data[1323] = ~16'b0;
    assign data[1324] = ~16'b0;
    assign data[1325] = ~16'b0;
    assign data[1326] = ~16'b0;
    assign data[1327] = ~16'b0;
    assign data[1328] = ~16'b0;
    assign data[1329] = ~16'b0;
    assign data[1330] = ~16'b0;
    assign data[1331] = ~16'b0;
    assign data[1332] = ~16'b0;
    assign data[1333] = ~16'b0;
    assign data[1334] = ~16'b0;
    assign data[1335] = ~16'b0;
    assign data[1336] = ~16'b0;
    assign data[1337] = ~16'b0;
    assign data[1338] = ~16'b0;
    assign data[1339] = ~16'b0;
    assign data[1340] = ~16'b0;
    assign data[1341] = ~16'b0;
    assign data[1342] = ~16'b0;
    assign data[1343] = ~16'b0;
    assign data[1344] = ~16'b0;
    assign data[1345] = ~16'b0;
    assign data[1346] = ~16'b0;
    assign data[1347] = ~16'b0;
    assign data[1348] = ~16'b0;
    assign data[1349] = ~16'b0;
    assign data[1350] = ~16'b0;
    assign data[1351] = ~16'b0;
    assign data[1352] = ~16'b0;
    assign data[1353] = ~16'b0;
    assign data[1354] = ~16'b0;
    assign data[1355] = ~16'b0;
    assign data[1356] = ~16'b0;
    assign data[1357] = ~16'b0;
    assign data[1358] = ~16'b0;
    assign data[1359] = ~16'b0;
    assign data[1360] = ~16'b0;
    assign data[1361] = ~16'b0;
    assign data[1362] = ~16'b0;
    assign data[1363] = ~16'b0;
    assign data[1364] = ~16'b0;
    assign data[1365] = ~16'b0;
    assign data[1366] = ~16'b0;
    assign data[1367] = ~16'b0;
    assign data[1368] = ~16'b0;
    assign data[1369] = ~16'b0;
    assign data[1370] = ~16'b0;
    assign data[1371] = ~16'b0;
    assign data[1372] = ~16'b0;
    assign data[1373] = ~16'b0;
    assign data[1374] = ~16'b0;
    assign data[1375] = ~16'b0;
    assign data[1376] = ~16'b0;
    assign data[1377] = ~16'b0;
    assign data[1378] = ~16'b0;
    assign data[1379] = ~16'b0;
    assign data[1380] = ~16'b0;
    assign data[1381] = ~16'b0;
    assign data[1382] = ~16'b0;
    assign data[1383] = ~16'b0;
    assign data[1384] = ~16'b0;
    assign data[1385] = ~16'b0;
    assign data[1386] = ~16'b0;
    assign data[1387] = ~16'b0;
    assign data[1388] = ~16'b0;
    assign data[1389] = ~16'b0;
    assign data[1390] = ~16'b0;
    assign data[1391] = ~16'b0;
    assign data[1392] = ~16'b0;
    assign data[1393] = ~16'b0;
    assign data[1394] = ~16'b0;
    assign data[1395] = ~16'b0;
    assign data[1396] = ~16'b0;
    assign data[1397] = ~16'b0;
    assign data[1398] = ~16'b0;
    assign data[1399] = ~16'b0;
    assign data[1400] = ~16'b0;
    assign data[1401] = ~16'b0;
    assign data[1402] = ~16'b0;
    assign data[1403] = ~16'b0;
    assign data[1404] = ~16'b0;
    assign data[1405] = ~16'b0;
    assign data[1406] = ~16'b0;
    assign data[1407] = ~16'b0;
    assign data[1408] = ~16'b0;
    assign data[1409] = ~16'b0;
    assign data[1410] = 16'b0;
    assign data[1411] = 16'b0;
    assign data[1412] = 16'b0;
    assign data[1413] = 16'b0;
    assign data[1414] = 16'b0;
    assign data[1415] = 16'b0;
    assign data[1416] = 16'b0;
    assign data[1417] = 16'b0;
    assign data[1418] = 16'b0;
    assign data[1419] = 16'b0;
    assign data[1420] = 16'b0;
    assign data[1421] = 16'b0;
    assign data[1422] = 16'b0;
    assign data[1423] = 16'b0;
    assign data[1424] = 16'b0;
    assign data[1425] = 16'b0;
    assign data[1426] = 16'b0;
    assign data[1427] = 16'b0;
    assign data[1428] = 16'b0;
    assign data[1429] = 16'b0;
    assign data[1430] = 16'b0;
    assign data[1431] = 16'b0;
    assign data[1432] = ~16'b0;
    assign data[1433] = ~16'b0;
    assign data[1434] = ~16'b0;
    assign data[1435] = ~16'b0;
    assign data[1436] = ~16'b0;
    assign data[1437] = ~16'b0;
    assign data[1438] = ~16'b0;
    assign data[1439] = ~16'b0;
    assign data[1440] = 16'b0;
    assign data[1441] = 16'b0;
    assign data[1442] = ~16'b0;
    assign data[1443] = ~16'b0;
    assign data[1444] = ~16'b0;
    assign data[1445] = ~16'b0;
    assign data[1446] = ~16'b0;
    assign data[1447] = ~16'b0;
    assign data[1448] = ~16'b0;
    assign data[1449] = ~16'b0;
    assign data[1450] = 16'b0;
    assign data[1451] = 16'b0;
    assign data[1452] = ~16'b0;
    assign data[1453] = ~16'b0;
    assign data[1454] = ~16'b0;
    assign data[1455] = ~16'b0;
    assign data[1456] = ~16'b0;
    assign data[1457] = ~16'b0;
    assign data[1458] = ~16'b0;
    assign data[1459] = ~16'b0;
    assign data[1460] = 16'b0;
    assign data[1461] = 16'b0;
    assign data[1462] = ~16'b0;
    assign data[1463] = ~16'b0;
    assign data[1464] = ~16'b0;
    assign data[1465] = ~16'b0;
    assign data[1466] = ~16'b0;
    assign data[1467] = ~16'b0;
    assign data[1468] = ~16'b0;
    assign data[1469] = ~16'b0;
    assign data[1470] = 16'b0;
    assign data[1471] = 16'b0;
    assign data[1472] = ~16'b0;
    assign data[1473] = ~16'b0;
    assign data[1474] = ~16'b0;
    assign data[1475] = ~16'b0;
    assign data[1476] = ~16'b0;
    assign data[1477] = ~16'b0;
    assign data[1478] = ~16'b0;
    assign data[1479] = ~16'b0;
    assign data[1480] = 16'b0;
    assign data[1481] = 16'b0;
    assign data[1482] = ~16'b0;
    assign data[1483] = ~16'b0;
    assign data[1484] = ~16'b0;
    assign data[1485] = ~16'b0;
    assign data[1486] = ~16'b0;
    assign data[1487] = ~16'b0;
    assign data[1488] = ~16'b0;
    assign data[1489] = ~16'b0;
    assign data[1490] = 16'b0;
    assign data[1491] = 16'b0;
    assign data[1492] = ~16'b0;
    assign data[1493] = ~16'b0;
    assign data[1494] = ~16'b0;
    assign data[1495] = ~16'b0;
    assign data[1496] = ~16'b0;
    assign data[1497] = ~16'b0;
    assign data[1498] = ~16'b0;
    assign data[1499] = ~16'b0;
    assign data[1500] = 16'b0;
    assign data[1501] = 16'b0;
    assign data[1502] = ~16'b0;
    assign data[1503] = ~16'b0;
    assign data[1504] = ~16'b0;
    assign data[1505] = ~16'b0;
    assign data[1506] = ~16'b0;
    assign data[1507] = ~16'b0;
    assign data[1508] = ~16'b0;
    assign data[1509] = ~16'b0;
    assign data[1510] = 16'b0;
    assign data[1511] = 16'b0;
    assign data[1512] = ~16'b0;
    assign data[1513] = ~16'b0;
    assign data[1514] = ~16'b0;
    assign data[1515] = ~16'b0;
    assign data[1516] = ~16'b0;
    assign data[1517] = ~16'b0;
    assign data[1518] = ~16'b0;
    assign data[1519] = ~16'b0;
    assign data[1520] = 16'b0;
    assign data[1521] = 16'b0;
    assign data[1522] = ~16'b0;
    assign data[1523] = ~16'b0;
    assign data[1524] = ~16'b0;
    assign data[1525] = ~16'b0;
    assign data[1526] = ~16'b0;
    assign data[1527] = ~16'b0;
    assign data[1528] = ~16'b0;
    assign data[1529] = ~16'b0;
    assign data[1530] = 16'b0;
    assign data[1531] = 16'b0;
    assign data[1532] = ~16'b0;
    assign data[1533] = ~16'b0;
    assign data[1534] = ~16'b0;
    assign data[1535] = ~16'b0;
    assign data[1536] = ~16'b0;
    assign data[1537] = ~16'b0;
    assign data[1538] = ~16'b0;
    assign data[1539] = ~16'b0;
    assign data[1540] = 16'b0;
    assign data[1541] = 16'b0;
    assign data[1542] = ~16'b0;
    assign data[1543] = ~16'b0;
    assign data[1544] = ~16'b0;
    assign data[1545] = ~16'b0;
    assign data[1546] = ~16'b0;
    assign data[1547] = ~16'b0;
    assign data[1548] = ~16'b0;
    assign data[1549] = ~16'b0;
    assign data[1550] = 16'b0;
    assign data[1551] = 16'b0;
    assign data[1552] = ~16'b0;
    assign data[1553] = ~16'b0;
    assign data[1554] = ~16'b0;
    assign data[1555] = ~16'b0;
    assign data[1556] = ~16'b0;
    assign data[1557] = ~16'b0;
    assign data[1558] = ~16'b0;
    assign data[1559] = ~16'b0;
    assign data[1560] = 16'b0;
    assign data[1561] = 16'b0;
    assign data[1562] = ~16'b0;
    assign data[1563] = ~16'b0;
    assign data[1564] = ~16'b0;
    assign data[1565] = ~16'b0;
    assign data[1566] = ~16'b0;
    assign data[1567] = ~16'b0;
    assign data[1568] = ~16'b0;
    assign data[1569] = ~16'b0;
    assign data[1570] = 16'b0;
    assign data[1571] = 16'b0;
    assign data[1572] = ~16'b0;
    assign data[1573] = ~16'b0;
    assign data[1574] = ~16'b0;
    assign data[1575] = ~16'b0;
    assign data[1576] = ~16'b0;
    assign data[1577] = ~16'b0;
    assign data[1578] = ~16'b0;
    assign data[1579] = ~16'b0;
    assign data[1580] = 16'b0;
    assign data[1581] = 16'b0;
    assign data[1582] = ~16'b0;
    assign data[1583] = ~16'b0;
    assign data[1584] = ~16'b0;
    assign data[1585] = ~16'b0;
    assign data[1586] = ~16'b0;
    assign data[1587] = ~16'b0;
    assign data[1588] = ~16'b0;
    assign data[1589] = ~16'b0;
    assign data[1590] = 16'b0;
    assign data[1591] = 16'b0;
    assign data[1592] = ~16'b0;
    assign data[1593] = ~16'b0;
    assign data[1594] = ~16'b0;
    assign data[1595] = ~16'b0;
    assign data[1596] = ~16'b0;
    assign data[1597] = ~16'b0;
    assign data[1598] = ~16'b0;
    assign data[1599] = ~16'b0;
    assign data[1600] = 16'b0;
    assign data[1601] = 16'b0;
    assign data[1602] = ~16'b0;
    assign data[1603] = ~16'b0;
    assign data[1604] = ~16'b0;
    assign data[1605] = ~16'b0;
    assign data[1606] = ~16'b0;
    assign data[1607] = ~16'b0;
    assign data[1608] = ~16'b0;
    assign data[1609] = ~16'b0;
    assign data[1610] = 16'b0;
    assign data[1611] = 16'b0;
    assign data[1612] = ~16'b0;
    assign data[1613] = ~16'b0;
    assign data[1614] = ~16'b0;
    assign data[1615] = ~16'b0;
    assign data[1616] = ~16'b0;
    assign data[1617] = ~16'b0;
    assign data[1618] = ~16'b0;
    assign data[1619] = ~16'b0;
    assign data[1620] = 16'b0;
    assign data[1621] = 16'b0;
    assign data[1622] = ~16'b0;
    assign data[1623] = ~16'b0;
    assign data[1624] = ~16'b0;
    assign data[1625] = ~16'b0;
    assign data[1626] = ~16'b0;
    assign data[1627] = ~16'b0;
    assign data[1628] = ~16'b0;
    assign data[1629] = ~16'b0;
    assign data[1630] = 16'b0;
    assign data[1631] = 16'b0;
    assign data[1632] = ~16'b0;
    assign data[1633] = ~16'b0;
    assign data[1634] = ~16'b0;
    assign data[1635] = ~16'b0;
    assign data[1636] = ~16'b0;
    assign data[1637] = ~16'b0;
    assign data[1638] = ~16'b0;
    assign data[1639] = ~16'b0;
    assign data[1640] = 16'b0;
    assign data[1641] = 16'b0;
    assign data[1642] = ~16'b0;
    assign data[1643] = ~16'b0;
    assign data[1644] = ~16'b0;
    assign data[1645] = ~16'b0;
    assign data[1646] = ~16'b0;
    assign data[1647] = ~16'b0;
    assign data[1648] = ~16'b0;
    assign data[1649] = ~16'b0;
    assign data[1650] = 16'b0;
    assign data[1651] = 16'b0;
    assign data[1652] = ~16'b0;
    assign data[1653] = ~16'b0;
    assign data[1654] = ~16'b0;
    assign data[1655] = ~16'b0;
    assign data[1656] = ~16'b0;
    assign data[1657] = ~16'b0;
    assign data[1658] = ~16'b0;
    assign data[1659] = ~16'b0;
    assign data[1660] = 16'b0;
    assign data[1661] = 16'b0;
    assign data[1662] = ~16'b0;
    assign data[1663] = ~16'b0;
    assign data[1664] = ~16'b0;
    assign data[1665] = ~16'b0;
    assign data[1666] = ~16'b0;
    assign data[1667] = ~16'b0;
    assign data[1668] = ~16'b0;
    assign data[1669] = ~16'b0;
    assign data[1670] = 16'b0;
    assign data[1671] = 16'b0;
    assign data[1672] = ~16'b0;
    assign data[1673] = ~16'b0;
    assign data[1674] = ~16'b0;
    assign data[1675] = ~16'b0;
    assign data[1676] = ~16'b0;
    assign data[1677] = ~16'b0;
    assign data[1678] = ~16'b0;
    assign data[1679] = ~16'b0;
    assign data[1680] = 16'b0;
    assign data[1681] = 16'b0;
    assign data[1682] = ~16'b0;
    assign data[1683] = ~16'b0;
    assign data[1684] = ~16'b0;
    assign data[1685] = ~16'b0;
    assign data[1686] = ~16'b0;
    assign data[1687] = ~16'b0;
    assign data[1688] = ~16'b0;
    assign data[1689] = ~16'b0;
    assign data[1690] = 16'b0;
    assign data[1691] = 16'b0;
    assign data[1692] = ~16'b0;
    assign data[1693] = ~16'b0;
    assign data[1694] = ~16'b0;
    assign data[1695] = ~16'b0;
    assign data[1696] = ~16'b0;
    assign data[1697] = ~16'b0;
    assign data[1698] = ~16'b0;
    assign data[1699] = ~16'b0;
    assign data[1700] = 16'b0;
    assign data[1701] = 16'b0;
    assign data[1702] = ~16'b0;
    assign data[1703] = ~16'b0;
    assign data[1704] = ~16'b0;
    assign data[1705] = ~16'b0;
    assign data[1706] = ~16'b0;
    assign data[1707] = ~16'b0;
    assign data[1708] = ~16'b0;
    assign data[1709] = ~16'b0;
    assign data[1710] = 16'b0;
    assign data[1711] = 16'b0;
    assign data[1712] = ~16'b0;
    assign data[1713] = ~16'b0;
    assign data[1714] = ~16'b0;
    assign data[1715] = ~16'b0;
    assign data[1716] = ~16'b0;
    assign data[1717] = ~16'b0;
    assign data[1718] = ~16'b0;
    assign data[1719] = ~16'b0;
    assign data[1720] = 16'b0;
    assign data[1721] = 16'b0;
    assign data[1722] = ~16'b0;
    assign data[1723] = ~16'b0;
    assign data[1724] = ~16'b0;
    assign data[1725] = ~16'b0;
    assign data[1726] = ~16'b0;
    assign data[1727] = ~16'b0;
    assign data[1728] = ~16'b0;
    assign data[1729] = ~16'b0;
    assign data[1730] = 16'b0;
    assign data[1731] = 16'b0;
    assign data[1732] = ~16'b0;
    assign data[1733] = ~16'b0;
    assign data[1734] = ~16'b0;
    assign data[1735] = ~16'b0;
    assign data[1736] = ~16'b0;
    assign data[1737] = ~16'b0;
    assign data[1738] = ~16'b0;
    assign data[1739] = ~16'b0;
    assign data[1740] = 16'b0;
    assign data[1741] = 16'b0;
    assign data[1742] = ~16'b0;
    assign data[1743] = ~16'b0;
    assign data[1744] = ~16'b0;
    assign data[1745] = ~16'b0;
    assign data[1746] = ~16'b0;
    assign data[1747] = ~16'b0;
    assign data[1748] = ~16'b0;
    assign data[1749] = ~16'b0;
    assign data[1750] = 16'b0;
    assign data[1751] = 16'b0;
    assign data[1752] = ~16'b0;
    assign data[1753] = ~16'b0;
    assign data[1754] = ~16'b0;
    assign data[1755] = ~16'b0;
    assign data[1756] = ~16'b0;
    assign data[1757] = ~16'b0;
    assign data[1758] = ~16'b0;
    assign data[1759] = ~16'b0;
    assign data[1760] = 16'b0;
    assign data[1761] = 16'b0;
    assign data[1762] = ~16'b0;
    assign data[1763] = ~16'b0;
    assign data[1764] = ~16'b0;
    assign data[1765] = ~16'b0;
    assign data[1766] = ~16'b0;
    assign data[1767] = ~16'b0;
    assign data[1768] = ~16'b0;
    assign data[1769] = ~16'b0;
    assign data[1770] = 16'b0;
    assign data[1771] = 16'b0;
    assign data[1772] = 16'b0;
    assign data[1773] = 16'b0;
    assign data[1774] = 16'b0;
    assign data[1775] = 16'b0;
    assign data[1776] = 16'b0;
    assign data[1777] = 16'b0;
    assign data[1778] = 16'b0;
    assign data[1779] = 16'b0;
    assign data[1780] = 16'b0;
    assign data[1781] = 16'b0;
    assign data[1782] = 16'b0;
    assign data[1783] = 16'b0;
    assign data[1784] = 16'b0;
    assign data[1785] = 16'b0;
    assign data[1786] = 16'b0;
    assign data[1787] = 16'b0;
    assign data[1788] = 16'b0;
    assign data[1789] = 16'b0;
    assign data[1790] = ~16'b0;
    assign data[1791] = ~16'b0;
    assign data[1792] = ~16'b0;
    assign data[1793] = ~16'b0;
    assign data[1794] = ~16'b0;
    assign data[1795] = ~16'b0;
    assign data[1796] = ~16'b0;
    assign data[1797] = ~16'b0;
    assign data[1798] = ~16'b0;
    assign data[1799] = ~16'b0;
    assign data[1800] = ~16'b0;
    assign data[1801] = ~16'b0;
    assign data[1802] = ~16'b0;
    assign data[1803] = ~16'b0;
    assign data[1804] = ~16'b0;
    assign data[1805] = ~16'b0;
    assign data[1806] = ~16'b0;
    assign data[1807] = ~16'b0;
    assign data[1808] = ~16'b0;
    assign data[1809] = ~16'b0;
    assign data[1810] = ~16'b0;
    assign data[1811] = ~16'b0;
    assign data[1812] = ~16'b0;
    assign data[1813] = ~16'b0;
    assign data[1814] = ~16'b0;
    assign data[1815] = ~16'b0;
    assign data[1816] = ~16'b0;
    assign data[1817] = ~16'b0;
    assign data[1818] = ~16'b0;
    assign data[1819] = ~16'b0;
    assign data[1820] = ~16'b0;
    assign data[1821] = ~16'b0;
    assign data[1822] = ~16'b0;
    assign data[1823] = ~16'b0;
    assign data[1824] = ~16'b0;
    assign data[1825] = ~16'b0;
    assign data[1826] = ~16'b0;
    assign data[1827] = ~16'b0;
    assign data[1828] = ~16'b0;
    assign data[1829] = ~16'b0;
    assign data[1830] = ~16'b0;
    assign data[1831] = ~16'b0;
    assign data[1832] = ~16'b0;
    assign data[1833] = ~16'b0;
    assign data[1834] = ~16'b0;
    assign data[1835] = ~16'b0;
    assign data[1836] = ~16'b0;
    assign data[1837] = ~16'b0;
    assign data[1838] = ~16'b0;
    assign data[1839] = ~16'b0;
    assign data[1840] = ~16'b0;
    assign data[1841] = ~16'b0;
    assign data[1842] = ~16'b0;
    assign data[1843] = ~16'b0;
    assign data[1844] = ~16'b0;
    assign data[1845] = ~16'b0;
    assign data[1846] = ~16'b0;
    assign data[1847] = ~16'b0;
    assign data[1848] = ~16'b0;
    assign data[1849] = ~16'b0;
    assign data[1850] = ~16'b0;
    assign data[1851] = ~16'b0;
    assign data[1852] = ~16'b0;
    assign data[1853] = ~16'b0;
    assign data[1854] = ~16'b0;
    assign data[1855] = ~16'b0;
    assign data[1856] = ~16'b0;
    assign data[1857] = ~16'b0;
    assign data[1858] = ~16'b0;
    assign data[1859] = ~16'b0;
    assign data[1860] = ~16'b0;
    assign data[1861] = ~16'b0;
    assign data[1862] = ~16'b0;
    assign data[1863] = ~16'b0;
    assign data[1864] = ~16'b0;
    assign data[1865] = ~16'b0;
    assign data[1866] = ~16'b0;
    assign data[1867] = ~16'b0;
    assign data[1868] = ~16'b0;
    assign data[1869] = ~16'b0;
    assign data[1870] = ~16'b0;
    assign data[1871] = ~16'b0;
    assign data[1872] = ~16'b0;
    assign data[1873] = ~16'b0;
    assign data[1874] = ~16'b0;
    assign data[1875] = ~16'b0;
    assign data[1876] = ~16'b0;
    assign data[1877] = ~16'b0;
    assign data[1878] = ~16'b0;
    assign data[1879] = ~16'b0;
    assign data[1880] = ~16'b0;
    assign data[1881] = ~16'b0;
    assign data[1882] = ~16'b0;
    assign data[1883] = ~16'b0;
    assign data[1884] = ~16'b0;
    assign data[1885] = ~16'b0;
    assign data[1886] = ~16'b0;
    assign data[1887] = ~16'b0;
    assign data[1888] = ~16'b0;
    assign data[1889] = ~16'b0;
    assign data[1890] = ~16'b0;
    assign data[1891] = ~16'b0;
    assign data[1892] = ~16'b0;
    assign data[1893] = ~16'b0;
    assign data[1894] = ~16'b0;
    assign data[1895] = ~16'b0;
    assign data[1896] = ~16'b0;
    assign data[1897] = ~16'b0;
    assign data[1898] = ~16'b0;
    assign data[1899] = ~16'b0;
    assign data[1900] = ~16'b0;
    assign data[1901] = ~16'b0;
    assign data[1902] = ~16'b0;
    assign data[1903] = ~16'b0;
    assign data[1904] = ~16'b0;
    assign data[1905] = ~16'b0;
    assign data[1906] = ~16'b0;
    assign data[1907] = ~16'b0;
    assign data[1908] = ~16'b0;
    assign data[1909] = ~16'b0;
    assign data[1910] = ~16'b0;
    assign data[1911] = ~16'b0;
    assign data[1912] = ~16'b0;
    assign data[1913] = ~16'b0;
    assign data[1914] = ~16'b0;
    assign data[1915] = ~16'b0;
    assign data[1916] = ~16'b0;
    assign data[1917] = ~16'b0;
    assign data[1918] = ~16'b0;
    assign data[1919] = ~16'b0;
    assign data[1920] = ~16'b0;
    assign data[1921] = ~16'b0;
    assign data[1922] = ~16'b0;
    assign data[1923] = ~16'b0;
    assign data[1924] = ~16'b0;
    assign data[1925] = ~16'b0;
    assign data[1926] = ~16'b0;
    assign data[1927] = ~16'b0;
    assign data[1928] = ~16'b0;
    assign data[1929] = ~16'b0;
    assign data[1930] = ~16'b0;
    assign data[1931] = ~16'b0;
    assign data[1932] = ~16'b0;
    assign data[1933] = ~16'b0;
    assign data[1934] = ~16'b0;
    assign data[1935] = ~16'b0;
    assign data[1936] = ~16'b0;
    assign data[1937] = ~16'b0;
    assign data[1938] = ~16'b0;
    assign data[1939] = ~16'b0;
    assign data[1940] = ~16'b0;
    assign data[1941] = ~16'b0;
    assign data[1942] = ~16'b0;
    assign data[1943] = ~16'b0;
    assign data[1944] = ~16'b0;
    assign data[1945] = ~16'b0;
    assign data[1946] = ~16'b0;
    assign data[1947] = ~16'b0;
    assign data[1948] = ~16'b0;
    assign data[1949] = ~16'b0;
    assign data[1950] = ~16'b0;
    assign data[1951] = ~16'b0;
    assign data[1952] = ~16'b0;
    assign data[1953] = ~16'b0;
    assign data[1954] = ~16'b0;
    assign data[1955] = ~16'b0;
    assign data[1956] = ~16'b0;
    assign data[1957] = ~16'b0;
    assign data[1958] = ~16'b0;
    assign data[1959] = ~16'b0;
    assign data[1960] = ~16'b0;
    assign data[1961] = ~16'b0;
    assign data[1962] = ~16'b0;
    assign data[1963] = ~16'b0;
    assign data[1964] = ~16'b0;
    assign data[1965] = ~16'b0;
    assign data[1966] = ~16'b0;
    assign data[1967] = ~16'b0;
    assign data[1968] = ~16'b0;
    assign data[1969] = ~16'b0;
    assign data[1970] = ~16'b0;
    assign data[1971] = ~16'b0;
    assign data[1972] = ~16'b0;
    assign data[1973] = ~16'b0;
    assign data[1974] = ~16'b0;
    assign data[1975] = ~16'b0;
    assign data[1976] = ~16'b0;
    assign data[1977] = ~16'b0;
    assign data[1978] = ~16'b0;
    assign data[1979] = ~16'b0;
    assign data[1980] = ~16'b0;
    assign data[1981] = ~16'b0;
    assign data[1982] = ~16'b0;
    assign data[1983] = ~16'b0;
    assign data[1984] = ~16'b0;
    assign data[1985] = ~16'b0;
    assign data[1986] = ~16'b0;
    assign data[1987] = ~16'b0;
    assign data[1988] = ~16'b0;
    assign data[1989] = ~16'b0;
    assign data[1990] = ~16'b0;
    assign data[1991] = ~16'b0;
    assign data[1992] = ~16'b0;
    assign data[1993] = ~16'b0;
    assign data[1994] = ~16'b0;
    assign data[1995] = ~16'b0;
    assign data[1996] = ~16'b0;
    assign data[1997] = ~16'b0;
    assign data[1998] = ~16'b0;
    assign data[1999] = ~16'b0;
    assign data[2000] = ~16'b0;
    assign data[2001] = ~16'b0;
    assign data[2002] = ~16'b0;
    assign data[2003] = ~16'b0;
    assign data[2004] = ~16'b0;
    assign data[2005] = ~16'b0;
    assign data[2006] = ~16'b0;
    assign data[2007] = ~16'b0;
    assign data[2008] = ~16'b0;
    assign data[2009] = ~16'b0;
    assign data[2010] = ~16'b0;
    assign data[2011] = ~16'b0;
    assign data[2012] = ~16'b0;
    assign data[2013] = ~16'b0;
    assign data[2014] = ~16'b0;
    assign data[2015] = ~16'b0;
    assign data[2016] = ~16'b0;
    assign data[2017] = ~16'b0;
    assign data[2018] = ~16'b0;
    assign data[2019] = ~16'b0;
    assign data[2020] = 16'b0;
    assign data[2021] = 16'b0;
    assign data[2022] = 16'b0;
    assign data[2023] = 16'b0;
    assign data[2024] = 16'b0;
    assign data[2025] = 16'b0;
    assign data[2026] = 16'b0;
    assign data[2027] = 16'b0;
    assign data[2028] = 16'b0;
    assign data[2029] = 16'b0;
    assign data[2030] = 16'b0;
    assign data[2031] = 16'b0;
    assign data[2032] = 16'b0;
    assign data[2033] = 16'b0;
    assign data[2034] = 16'b0;
    assign data[2035] = 16'b0;
    assign data[2036] = 16'b0;
    assign data[2037] = 16'b0;
    assign data[2038] = 16'b0;
    assign data[2039] = 16'b0;
    assign data[2040] = 16'b0;
    assign data[2041] = 16'b0;
    assign data[2042] = ~16'b0;
    assign data[2043] = ~16'b0;
    assign data[2044] = ~16'b0;
    assign data[2045] = ~16'b0;
    assign data[2046] = ~16'b0;
    assign data[2047] = ~16'b0;
    assign data[2048] = ~16'b0;
    assign data[2049] = ~16'b0;
    assign data[2050] = 16'b0;
    assign data[2051] = 16'b0;
    assign data[2052] = ~16'b0;
    assign data[2053] = ~16'b0;
    assign data[2054] = ~16'b0;
    assign data[2055] = ~16'b0;
    assign data[2056] = ~16'b0;
    assign data[2057] = ~16'b0;
    assign data[2058] = ~16'b0;
    assign data[2059] = ~16'b0;
    assign data[2060] = 16'b0;
    assign data[2061] = 16'b0;
    assign data[2062] = ~16'b0;
    assign data[2063] = ~16'b0;
    assign data[2064] = ~16'b0;
    assign data[2065] = ~16'b0;
    assign data[2066] = ~16'b0;
    assign data[2067] = ~16'b0;
    assign data[2068] = ~16'b0;
    assign data[2069] = ~16'b0;
    assign data[2070] = 16'b0;
    assign data[2071] = 16'b0;
    assign data[2072] = ~16'b0;
    assign data[2073] = ~16'b0;
    assign data[2074] = ~16'b0;
    assign data[2075] = ~16'b0;
    assign data[2076] = ~16'b0;
    assign data[2077] = ~16'b0;
    assign data[2078] = ~16'b0;
    assign data[2079] = ~16'b0;
    assign data[2080] = 16'b0;
    assign data[2081] = 16'b0;
    assign data[2082] = ~16'b0;
    assign data[2083] = ~16'b0;
    assign data[2084] = ~16'b0;
    assign data[2085] = ~16'b0;
    assign data[2086] = ~16'b0;
    assign data[2087] = ~16'b0;
    assign data[2088] = ~16'b0;
    assign data[2089] = ~16'b0;
    assign data[2090] = 16'b0;
    assign data[2091] = 16'b0;
    assign data[2092] = ~16'b0;
    assign data[2093] = ~16'b0;
    assign data[2094] = ~16'b0;
    assign data[2095] = ~16'b0;
    assign data[2096] = ~16'b0;
    assign data[2097] = ~16'b0;
    assign data[2098] = ~16'b0;
    assign data[2099] = ~16'b0;
    assign data[2100] = 16'b0;
    assign data[2101] = 16'b0;
    assign data[2102] = ~16'b0;
    assign data[2103] = ~16'b0;
    assign data[2104] = ~16'b0;
    assign data[2105] = ~16'b0;
    assign data[2106] = ~16'b0;
    assign data[2107] = ~16'b0;
    assign data[2108] = ~16'b0;
    assign data[2109] = ~16'b0;
    assign data[2110] = 16'b0;
    assign data[2111] = 16'b0;
    assign data[2112] = ~16'b0;
    assign data[2113] = ~16'b0;
    assign data[2114] = ~16'b0;
    assign data[2115] = ~16'b0;
    assign data[2116] = ~16'b0;
    assign data[2117] = ~16'b0;
    assign data[2118] = ~16'b0;
    assign data[2119] = ~16'b0;
    assign data[2120] = 16'b0;
    assign data[2121] = 16'b0;
    assign data[2122] = ~16'b0;
    assign data[2123] = ~16'b0;
    assign data[2124] = ~16'b0;
    assign data[2125] = ~16'b0;
    assign data[2126] = ~16'b0;
    assign data[2127] = ~16'b0;
    assign data[2128] = ~16'b0;
    assign data[2129] = ~16'b0;
    assign data[2130] = 16'b0;
    assign data[2131] = 16'b0;
    assign data[2132] = ~16'b0;
    assign data[2133] = ~16'b0;
    assign data[2134] = ~16'b0;
    assign data[2135] = ~16'b0;
    assign data[2136] = ~16'b0;
    assign data[2137] = ~16'b0;
    assign data[2138] = ~16'b0;
    assign data[2139] = ~16'b0;
    assign data[2140] = 16'b0;
    assign data[2141] = 16'b0;
    assign data[2142] = ~16'b0;
    assign data[2143] = ~16'b0;
    assign data[2144] = ~16'b0;
    assign data[2145] = ~16'b0;
    assign data[2146] = ~16'b0;
    assign data[2147] = ~16'b0;
    assign data[2148] = ~16'b0;
    assign data[2149] = ~16'b0;
    assign data[2150] = 16'b0;
    assign data[2151] = 16'b0;
    assign data[2152] = ~16'b0;
    assign data[2153] = ~16'b0;
    assign data[2154] = ~16'b0;
    assign data[2155] = ~16'b0;
    assign data[2156] = ~16'b0;
    assign data[2157] = ~16'b0;
    assign data[2158] = ~16'b0;
    assign data[2159] = ~16'b0;
    assign data[2160] = 16'b0;
    assign data[2161] = 16'b0;
    assign data[2162] = ~16'b0;
    assign data[2163] = ~16'b0;
    assign data[2164] = ~16'b0;
    assign data[2165] = ~16'b0;
    assign data[2166] = ~16'b0;
    assign data[2167] = ~16'b0;
    assign data[2168] = ~16'b0;
    assign data[2169] = ~16'b0;
    assign data[2170] = 16'b0;
    assign data[2171] = 16'b0;
    assign data[2172] = ~16'b0;
    assign data[2173] = ~16'b0;
    assign data[2174] = ~16'b0;
    assign data[2175] = ~16'b0;
    assign data[2176] = ~16'b0;
    assign data[2177] = ~16'b0;
    assign data[2178] = ~16'b0;
    assign data[2179] = ~16'b0;
    assign data[2180] = 16'b0;
    assign data[2181] = 16'b0;
    assign data[2182] = ~16'b0;
    assign data[2183] = ~16'b0;
    assign data[2184] = ~16'b0;
    assign data[2185] = ~16'b0;
    assign data[2186] = ~16'b0;
    assign data[2187] = ~16'b0;
    assign data[2188] = ~16'b0;
    assign data[2189] = ~16'b0;
    assign data[2190] = 16'b0;
    assign data[2191] = 16'b0;
    assign data[2192] = ~16'b0;
    assign data[2193] = ~16'b0;
    assign data[2194] = ~16'b0;
    assign data[2195] = ~16'b0;
    assign data[2196] = ~16'b0;
    assign data[2197] = ~16'b0;
    assign data[2198] = ~16'b0;
    assign data[2199] = ~16'b0;
    assign data[2200] = 16'b0;
    assign data[2201] = 16'b0;
    assign data[2202] = 16'b0;
    assign data[2203] = 16'b0;
    assign data[2204] = 16'b0;
    assign data[2205] = 16'b0;
    assign data[2206] = 16'b0;
    assign data[2207] = 16'b0;
    assign data[2208] = 16'b0;
    assign data[2209] = 16'b0;
    assign data[2210] = 16'b0;
    assign data[2211] = 16'b0;
    assign data[2212] = 16'b0;
    assign data[2213] = 16'b0;
    assign data[2214] = 16'b0;
    assign data[2215] = 16'b0;
    assign data[2216] = 16'b0;
    assign data[2217] = 16'b0;
    assign data[2218] = 16'b0;
    assign data[2219] = 16'b0;
    assign data[2220] = ~16'b0;
    assign data[2221] = ~16'b0;
    assign data[2222] = ~16'b0;
    assign data[2223] = ~16'b0;
    assign data[2224] = ~16'b0;
    assign data[2225] = ~16'b0;
    assign data[2226] = ~16'b0;
    assign data[2227] = ~16'b0;
    assign data[2228] = ~16'b0;
    assign data[2229] = ~16'b0;
    assign data[2230] = ~16'b0;
    assign data[2231] = ~16'b0;
    assign data[2232] = ~16'b0;
    assign data[2233] = ~16'b0;
    assign data[2234] = ~16'b0;
    assign data[2235] = ~16'b0;
    assign data[2236] = ~16'b0;
    assign data[2237] = ~16'b0;
    assign data[2238] = ~16'b0;
    assign data[2239] = ~16'b0;
    assign data[2240] = ~16'b0;
    assign data[2241] = ~16'b0;
    assign data[2242] = ~16'b0;
    assign data[2243] = ~16'b0;
    assign data[2244] = ~16'b0;
    assign data[2245] = ~16'b0;
    assign data[2246] = ~16'b0;
    assign data[2247] = ~16'b0;
    assign data[2248] = ~16'b0;
    assign data[2249] = ~16'b0;
    assign data[2250] = ~16'b0;
    assign data[2251] = ~16'b0;
    assign data[2252] = ~16'b0;
    assign data[2253] = ~16'b0;
    assign data[2254] = ~16'b0;
    assign data[2255] = ~16'b0;
    assign data[2256] = ~16'b0;
    assign data[2257] = ~16'b0;
    assign data[2258] = ~16'b0;
    assign data[2259] = ~16'b0;
    assign data[2260] = ~16'b0;
    assign data[2261] = ~16'b0;
    assign data[2262] = ~16'b0;
    assign data[2263] = ~16'b0;
    assign data[2264] = ~16'b0;
    assign data[2265] = ~16'b0;
    assign data[2266] = ~16'b0;
    assign data[2267] = ~16'b0;
    assign data[2268] = ~16'b0;
    assign data[2269] = ~16'b0;
    assign data[2270] = ~16'b0;
    assign data[2271] = ~16'b0;
    assign data[2272] = ~16'b0;
    assign data[2273] = ~16'b0;
    assign data[2274] = ~16'b0;
    assign data[2275] = ~16'b0;
    assign data[2276] = ~16'b0;
    assign data[2277] = ~16'b0;
    assign data[2278] = ~16'b0;
    assign data[2279] = ~16'b0;
    assign data[2280] = ~16'b0;
    assign data[2281] = ~16'b0;
    assign data[2282] = ~16'b0;
    assign data[2283] = ~16'b0;
    assign data[2284] = ~16'b0;
    assign data[2285] = ~16'b0;
    assign data[2286] = ~16'b0;
    assign data[2287] = ~16'b0;
    assign data[2288] = ~16'b0;
    assign data[2289] = ~16'b0;
    assign data[2290] = ~16'b0;
    assign data[2291] = ~16'b0;
    assign data[2292] = ~16'b0;
    assign data[2293] = ~16'b0;
    assign data[2294] = ~16'b0;
    assign data[2295] = ~16'b0;
    assign data[2296] = ~16'b0;
    assign data[2297] = ~16'b0;
    assign data[2298] = ~16'b0;
    assign data[2299] = ~16'b0;
    assign data[2300] = ~16'b0;
    assign data[2301] = ~16'b0;
    assign data[2302] = ~16'b0;
    assign data[2303] = ~16'b0;
    assign data[2304] = ~16'b0;
    assign data[2305] = ~16'b0;
    assign data[2306] = ~16'b0;
    assign data[2307] = ~16'b0;
    assign data[2308] = ~16'b0;
    assign data[2309] = ~16'b0;
    assign data[2310] = ~16'b0;
    assign data[2311] = ~16'b0;
    assign data[2312] = ~16'b0;
    assign data[2313] = ~16'b0;
    assign data[2314] = ~16'b0;
    assign data[2315] = ~16'b0;
    assign data[2316] = ~16'b0;
    assign data[2317] = ~16'b0;
    assign data[2318] = ~16'b0;
    assign data[2319] = ~16'b0;
    assign data[2320] = 16'b0;
    assign data[2321] = 16'b0;
    assign data[2322] = 16'b0;
    assign data[2323] = 16'b0;
    assign data[2324] = 16'b0;
    assign data[2325] = 16'b0;
    assign data[2326] = 16'b0;
    assign data[2327] = 16'b0;
    assign data[2328] = 16'b0;
    assign data[2329] = 16'b0;
    assign data[2330] = 16'b0;
    assign data[2331] = 16'b0;
    assign data[2332] = 16'b0;
    assign data[2333] = 16'b0;
    assign data[2334] = 16'b0;
    assign data[2335] = 16'b0;
    assign data[2336] = 16'b0;
    assign data[2337] = 16'b0;
    assign data[2338] = 16'b0;
    assign data[2339] = 16'b0;
    assign data[2340] = 16'b0;
    assign data[2341] = 16'b0;
    assign data[2342] = ~16'b0;
    assign data[2343] = ~16'b0;
    assign data[2344] = ~16'b0;
    assign data[2345] = ~16'b0;
    assign data[2346] = ~16'b0;
    assign data[2347] = ~16'b0;
    assign data[2348] = ~16'b0;
    assign data[2349] = ~16'b0;
    assign data[2350] = 16'b0;
    assign data[2351] = 16'b0;
    assign data[2352] = ~16'b0;
    assign data[2353] = ~16'b0;
    assign data[2354] = ~16'b0;
    assign data[2355] = ~16'b0;
    assign data[2356] = ~16'b0;
    assign data[2357] = ~16'b0;
    assign data[2358] = ~16'b0;
    assign data[2359] = ~16'b0;
    assign data[2360] = 16'b0;
    assign data[2361] = 16'b0;
    assign data[2362] = ~16'b0;
    assign data[2363] = ~16'b0;
    assign data[2364] = ~16'b0;
    assign data[2365] = ~16'b0;
    assign data[2366] = ~16'b0;
    assign data[2367] = ~16'b0;
    assign data[2368] = ~16'b0;
    assign data[2369] = ~16'b0;
    assign data[2370] = 16'b0;
    assign data[2371] = 16'b0;
    assign data[2372] = ~16'b0;
    assign data[2373] = ~16'b0;
    assign data[2374] = ~16'b0;
    assign data[2375] = ~16'b0;
    assign data[2376] = ~16'b0;
    assign data[2377] = ~16'b0;
    assign data[2378] = ~16'b0;
    assign data[2379] = ~16'b0;
    assign data[2380] = 16'b0;
    assign data[2381] = 16'b0;
    assign data[2382] = ~16'b0;
    assign data[2383] = ~16'b0;
    assign data[2384] = ~16'b0;
    assign data[2385] = ~16'b0;
    assign data[2386] = ~16'b0;
    assign data[2387] = ~16'b0;
    assign data[2388] = ~16'b0;
    assign data[2389] = ~16'b0;
    assign data[2390] = 16'b0;
    assign data[2391] = 16'b0;
    assign data[2392] = ~16'b0;
    assign data[2393] = ~16'b0;
    assign data[2394] = ~16'b0;
    assign data[2395] = ~16'b0;
    assign data[2396] = ~16'b0;
    assign data[2397] = ~16'b0;
    assign data[2398] = ~16'b0;
    assign data[2399] = ~16'b0;
    assign data[2400] = 16'b0;
    assign data[2401] = 16'b0;
    assign data[2402] = ~16'b0;
    assign data[2403] = ~16'b0;
    assign data[2404] = ~16'b0;
    assign data[2405] = ~16'b0;
    assign data[2406] = ~16'b0;
    assign data[2407] = ~16'b0;
    assign data[2408] = ~16'b0;
    assign data[2409] = ~16'b0;
    assign data[2410] = 16'b0;
    assign data[2411] = 16'b0;
    assign data[2412] = ~16'b0;
    assign data[2413] = ~16'b0;
    assign data[2414] = ~16'b0;
    assign data[2415] = ~16'b0;
    assign data[2416] = ~16'b0;
    assign data[2417] = ~16'b0;
    assign data[2418] = ~16'b0;
    assign data[2419] = ~16'b0;
    assign data[2420] = 16'b0;
    assign data[2421] = 16'b0;
    assign data[2422] = ~16'b0;
    assign data[2423] = ~16'b0;
    assign data[2424] = ~16'b0;
    assign data[2425] = ~16'b0;
    assign data[2426] = ~16'b0;
    assign data[2427] = ~16'b0;
    assign data[2428] = ~16'b0;
    assign data[2429] = ~16'b0;
    assign data[2430] = 16'b0;
    assign data[2431] = 16'b0;
    assign data[2432] = ~16'b0;
    assign data[2433] = ~16'b0;
    assign data[2434] = ~16'b0;
    assign data[2435] = ~16'b0;
    assign data[2436] = ~16'b0;
    assign data[2437] = ~16'b0;
    assign data[2438] = ~16'b0;
    assign data[2439] = ~16'b0;
    assign data[2440] = 16'b0;
    assign data[2441] = 16'b0;
    assign data[2442] = ~16'b0;
    assign data[2443] = ~16'b0;
    assign data[2444] = ~16'b0;
    assign data[2445] = ~16'b0;
    assign data[2446] = ~16'b0;
    assign data[2447] = ~16'b0;
    assign data[2448] = ~16'b0;
    assign data[2449] = ~16'b0;
    assign data[2450] = 16'b0;
    assign data[2451] = 16'b0;
    assign data[2452] = ~16'b0;
    assign data[2453] = ~16'b0;
    assign data[2454] = ~16'b0;
    assign data[2455] = ~16'b0;
    assign data[2456] = ~16'b0;
    assign data[2457] = ~16'b0;
    assign data[2458] = ~16'b0;
    assign data[2459] = ~16'b0;
    assign data[2460] = 16'b0;
    assign data[2461] = 16'b0;
    assign data[2462] = ~16'b0;
    assign data[2463] = ~16'b0;
    assign data[2464] = ~16'b0;
    assign data[2465] = ~16'b0;
    assign data[2466] = ~16'b0;
    assign data[2467] = ~16'b0;
    assign data[2468] = ~16'b0;
    assign data[2469] = ~16'b0;
    assign data[2470] = 16'b0;
    assign data[2471] = 16'b0;
    assign data[2472] = ~16'b0;
    assign data[2473] = ~16'b0;
    assign data[2474] = ~16'b0;
    assign data[2475] = ~16'b0;
    assign data[2476] = ~16'b0;
    assign data[2477] = ~16'b0;
    assign data[2478] = ~16'b0;
    assign data[2479] = ~16'b0;
    assign data[2480] = 16'b0;
    assign data[2481] = 16'b0;
    assign data[2482] = ~16'b0;
    assign data[2483] = ~16'b0;
    assign data[2484] = ~16'b0;
    assign data[2485] = ~16'b0;
    assign data[2486] = ~16'b0;
    assign data[2487] = ~16'b0;
    assign data[2488] = ~16'b0;
    assign data[2489] = ~16'b0;
    assign data[2490] = 16'b0;
    assign data[2491] = 16'b0;
    assign data[2492] = ~16'b0;
    assign data[2493] = ~16'b0;
    assign data[2494] = ~16'b0;
    assign data[2495] = ~16'b0;
    assign data[2496] = ~16'b0;
    assign data[2497] = ~16'b0;
    assign data[2498] = ~16'b0;
    assign data[2499] = ~16'b0;
    assign data[2500] = 16'b0;
    assign data[2501] = 16'b0;
    assign data[2502] = ~16'b0;
    assign data[2503] = ~16'b0;
    assign data[2504] = ~16'b0;
    assign data[2505] = ~16'b0;
    assign data[2506] = ~16'b0;
    assign data[2507] = ~16'b0;
    assign data[2508] = ~16'b0;
    assign data[2509] = ~16'b0;
    assign data[2510] = 16'b0;
    assign data[2511] = 16'b0;
    assign data[2512] = 16'b0;
    assign data[2513] = 16'b0;
    assign data[2514] = 16'b0;
    assign data[2515] = 16'b0;
    assign data[2516] = 16'b0;
    assign data[2517] = 16'b0;
    assign data[2518] = 16'b0;
    assign data[2519] = 16'b0;
    assign data[2520] = 16'b0;
    assign data[2521] = 16'b0;
    assign data[2522] = 16'b0;
    assign data[2523] = 16'b0;
    assign data[2524] = 16'b0;
    assign data[2525] = 16'b0;
    assign data[2526] = 16'b0;
    assign data[2527] = 16'b0;
    assign data[2528] = 16'b0;
    assign data[2529] = 16'b0;
    assign data[2530] = ~16'b0;
    assign data[2531] = ~16'b0;
    assign data[2532] = ~16'b0;
    assign data[2533] = ~16'b0;
    assign data[2534] = ~16'b0;
    assign data[2535] = ~16'b0;
    assign data[2536] = ~16'b0;
    assign data[2537] = ~16'b0;
    assign data[2538] = ~16'b0;
    assign data[2539] = ~16'b0;
    assign data[2540] = ~16'b0;
    assign data[2541] = ~16'b0;
    assign data[2542] = ~16'b0;
    assign data[2543] = ~16'b0;
    assign data[2544] = ~16'b0;
    assign data[2545] = ~16'b0;
    assign data[2546] = ~16'b0;
    assign data[2547] = ~16'b0;
    assign data[2548] = ~16'b0;
    assign data[2549] = ~16'b0;
    assign data[2550] = ~16'b0;
    assign data[2551] = ~16'b0;
    assign data[2552] = ~16'b0;
    assign data[2553] = ~16'b0;
    assign data[2554] = ~16'b0;
    assign data[2555] = ~16'b0;
    assign data[2556] = ~16'b0;
    assign data[2557] = ~16'b0;
    assign data[2558] = ~16'b0;
    assign data[2559] = ~16'b0;
    assign data[2560] = ~16'b0;
    assign data[2561] = ~16'b0;
    assign data[2562] = ~16'b0;
    assign data[2563] = ~16'b0;
    assign data[2564] = ~16'b0;
    assign data[2565] = ~16'b0;
    assign data[2566] = ~16'b0;
    assign data[2567] = ~16'b0;
    assign data[2568] = ~16'b0;
    assign data[2569] = ~16'b0;
    assign data[2570] = ~16'b0;
    assign data[2571] = ~16'b0;
    assign data[2572] = ~16'b0;
    assign data[2573] = ~16'b0;
    assign data[2574] = ~16'b0;
    assign data[2575] = ~16'b0;
    assign data[2576] = ~16'b0;
    assign data[2577] = ~16'b0;
    assign data[2578] = ~16'b0;
    assign data[2579] = ~16'b0;
    assign data[2580] = ~16'b0;
    assign data[2581] = ~16'b0;
    assign data[2582] = ~16'b0;
    assign data[2583] = ~16'b0;
    assign data[2584] = ~16'b0;
    assign data[2585] = ~16'b0;
    assign data[2586] = ~16'b0;
    assign data[2587] = ~16'b0;
    assign data[2588] = ~16'b0;
    assign data[2589] = ~16'b0;
    assign data[2590] = ~16'b0;
    assign data[2591] = ~16'b0;
    assign data[2592] = ~16'b0;
    assign data[2593] = ~16'b0;
    assign data[2594] = ~16'b0;
    assign data[2595] = ~16'b0;
    assign data[2596] = ~16'b0;
    assign data[2597] = ~16'b0;
    assign data[2598] = ~16'b0;
    assign data[2599] = ~16'b0;
    assign data[2600] = ~16'b0;
    assign data[2601] = ~16'b0;
    assign data[2602] = ~16'b0;
    assign data[2603] = ~16'b0;
    assign data[2604] = ~16'b0;
    assign data[2605] = ~16'b0;
    assign data[2606] = ~16'b0;
    assign data[2607] = ~16'b0;
    assign data[2608] = ~16'b0;
    assign data[2609] = ~16'b0;
    assign data[2610] = ~16'b0;
    assign data[2611] = ~16'b0;
    assign data[2612] = ~16'b0;
    assign data[2613] = ~16'b0;
    assign data[2614] = ~16'b0;
    assign data[2615] = ~16'b0;
    assign data[2616] = ~16'b0;
    assign data[2617] = ~16'b0;
    assign data[2618] = ~16'b0;
    assign data[2619] = ~16'b0;
    assign data[2620] = ~16'b0;
    assign data[2621] = ~16'b0;
    assign data[2622] = ~16'b0;
    assign data[2623] = ~16'b0;
    assign data[2624] = ~16'b0;
    assign data[2625] = ~16'b0;
    assign data[2626] = ~16'b0;
    assign data[2627] = ~16'b0;
    assign data[2628] = ~16'b0;
    assign data[2629] = ~16'b0;
    assign data[2630] = ~16'b0;
    assign data[2631] = ~16'b0;
    assign data[2632] = ~16'b0;
    assign data[2633] = ~16'b0;
    assign data[2634] = ~16'b0;
    assign data[2635] = ~16'b0;
    assign data[2636] = ~16'b0;
    assign data[2637] = ~16'b0;
    assign data[2638] = ~16'b0;
    assign data[2639] = ~16'b0;
    assign data[2640] = ~16'b0;
    assign data[2641] = ~16'b0;
    assign data[2642] = ~16'b0;
    assign data[2643] = ~16'b0;
    assign data[2644] = ~16'b0;
    assign data[2645] = ~16'b0;
    assign data[2646] = ~16'b0;
    assign data[2647] = ~16'b0;
    assign data[2648] = ~16'b0;
    assign data[2649] = ~16'b0;
    assign data[2650] = ~16'b0;
    assign data[2651] = ~16'b0;
    assign data[2652] = ~16'b0;
    assign data[2653] = ~16'b0;
    assign data[2654] = ~16'b0;
    assign data[2655] = ~16'b0;
    assign data[2656] = ~16'b0;
    assign data[2657] = ~16'b0;
    assign data[2658] = ~16'b0;
    assign data[2659] = ~16'b0;
    assign data[2660] = ~16'b0;
    assign data[2661] = ~16'b0;
    assign data[2662] = ~16'b0;
    assign data[2663] = ~16'b0;
    assign data[2664] = ~16'b0;
    assign data[2665] = ~16'b0;
    assign data[2666] = ~16'b0;
    assign data[2667] = ~16'b0;
    assign data[2668] = ~16'b0;
    assign data[2669] = ~16'b0;
    assign data[2670] = ~16'b0;
    assign data[2671] = ~16'b0;
    assign data[2672] = ~16'b0;
    assign data[2673] = ~16'b0;
    assign data[2674] = ~16'b0;
    assign data[2675] = ~16'b0;
    assign data[2676] = ~16'b0;
    assign data[2677] = ~16'b0;
    assign data[2678] = ~16'b0;
    assign data[2679] = ~16'b0;
    assign data[2680] = ~16'b0;
    assign data[2681] = ~16'b0;
    assign data[2682] = ~16'b0;
    assign data[2683] = ~16'b0;
    assign data[2684] = ~16'b0;
    assign data[2685] = ~16'b0;
    assign data[2686] = ~16'b0;
    assign data[2687] = ~16'b0;
    assign data[2688] = ~16'b0;
    assign data[2689] = ~16'b0;
    assign data[2690] = ~16'b0;
    assign data[2691] = ~16'b0;
    assign data[2692] = ~16'b0;
    assign data[2693] = ~16'b0;
    assign data[2694] = ~16'b0;
    assign data[2695] = ~16'b0;
    assign data[2696] = ~16'b0;
    assign data[2697] = ~16'b0;
    assign data[2698] = ~16'b0;
    assign data[2699] = ~16'b0;
    assign data[2700] = 16'b0;
    assign data[2701] = 16'b0;
    assign data[2702] = 16'b0;
    assign data[2703] = 16'b0;
    assign data[2704] = 16'b0;
    assign data[2705] = 16'b0;
    assign data[2706] = 16'b0;
    assign data[2707] = 16'b0;
    assign data[2708] = 16'b0;
    assign data[2709] = 16'b0;
    assign data[2710] = 16'b0;
    assign data[2711] = 16'b0;
    assign data[2712] = 16'b0;
    assign data[2713] = 16'b0;
    assign data[2714] = 16'b0;
    assign data[2715] = 16'b0;
    assign data[2716] = 16'b0;
    assign data[2717] = 16'b0;
    assign data[2718] = 16'b0;
    assign data[2719] = 16'b0;
    assign data[2720] = 16'b0;
    assign data[2721] = 16'b0;
    assign data[2722] = ~16'b0;
    assign data[2723] = ~16'b0;
    assign data[2724] = ~16'b0;
    assign data[2725] = ~16'b0;
    assign data[2726] = ~16'b0;
    assign data[2727] = ~16'b0;
    assign data[2728] = ~16'b0;
    assign data[2729] = ~16'b0;
    assign data[2730] = 16'b0;
    assign data[2731] = 16'b0;
    assign data[2732] = ~16'b0;
    assign data[2733] = ~16'b0;
    assign data[2734] = ~16'b0;
    assign data[2735] = ~16'b0;
    assign data[2736] = ~16'b0;
    assign data[2737] = ~16'b0;
    assign data[2738] = ~16'b0;
    assign data[2739] = ~16'b0;
    assign data[2740] = 16'b0;
    assign data[2741] = 16'b0;
    assign data[2742] = ~16'b0;
    assign data[2743] = ~16'b0;
    assign data[2744] = ~16'b0;
    assign data[2745] = ~16'b0;
    assign data[2746] = ~16'b0;
    assign data[2747] = ~16'b0;
    assign data[2748] = ~16'b0;
    assign data[2749] = ~16'b0;
    assign data[2750] = 16'b0;
    assign data[2751] = 16'b0;
    assign data[2752] = ~16'b0;
    assign data[2753] = ~16'b0;
    assign data[2754] = ~16'b0;
    assign data[2755] = ~16'b0;
    assign data[2756] = ~16'b0;
    assign data[2757] = ~16'b0;
    assign data[2758] = ~16'b0;
    assign data[2759] = ~16'b0;
    assign data[2760] = 16'b0;
    assign data[2761] = 16'b0;
    assign data[2762] = ~16'b0;
    assign data[2763] = ~16'b0;
    assign data[2764] = ~16'b0;
    assign data[2765] = ~16'b0;
    assign data[2766] = ~16'b0;
    assign data[2767] = ~16'b0;
    assign data[2768] = ~16'b0;
    assign data[2769] = ~16'b0;
    assign data[2770] = 16'b0;
    assign data[2771] = 16'b0;
    assign data[2772] = ~16'b0;
    assign data[2773] = ~16'b0;
    assign data[2774] = ~16'b0;
    assign data[2775] = ~16'b0;
    assign data[2776] = ~16'b0;
    assign data[2777] = ~16'b0;
    assign data[2778] = ~16'b0;
    assign data[2779] = ~16'b0;
    assign data[2780] = 16'b0;
    assign data[2781] = 16'b0;
    assign data[2782] = ~16'b0;
    assign data[2783] = ~16'b0;
    assign data[2784] = ~16'b0;
    assign data[2785] = ~16'b0;
    assign data[2786] = ~16'b0;
    assign data[2787] = ~16'b0;
    assign data[2788] = ~16'b0;
    assign data[2789] = ~16'b0;
    assign data[2790] = 16'b0;
    assign data[2791] = 16'b0;
    assign data[2792] = ~16'b0;
    assign data[2793] = ~16'b0;
    assign data[2794] = ~16'b0;
    assign data[2795] = ~16'b0;
    assign data[2796] = ~16'b0;
    assign data[2797] = ~16'b0;
    assign data[2798] = ~16'b0;
    assign data[2799] = ~16'b0;
    assign data[2800] = 16'b0;
    assign data[2801] = 16'b0;
    assign data[2802] = ~16'b0;
    assign data[2803] = ~16'b0;
    assign data[2804] = ~16'b0;
    assign data[2805] = ~16'b0;
    assign data[2806] = ~16'b0;
    assign data[2807] = ~16'b0;
    assign data[2808] = ~16'b0;
    assign data[2809] = ~16'b0;
    assign data[2810] = 16'b0;
    assign data[2811] = 16'b0;
    assign data[2812] = ~16'b0;
    assign data[2813] = ~16'b0;
    assign data[2814] = ~16'b0;
    assign data[2815] = ~16'b0;
    assign data[2816] = ~16'b0;
    assign data[2817] = ~16'b0;
    assign data[2818] = ~16'b0;
    assign data[2819] = ~16'b0;
    assign data[2820] = 16'b0;
    assign data[2821] = 16'b0;
    assign data[2822] = ~16'b0;
    assign data[2823] = ~16'b0;
    assign data[2824] = ~16'b0;
    assign data[2825] = ~16'b0;
    assign data[2826] = ~16'b0;
    assign data[2827] = ~16'b0;
    assign data[2828] = ~16'b0;
    assign data[2829] = ~16'b0;
    assign data[2830] = 16'b0;
    assign data[2831] = 16'b0;
    assign data[2832] = ~16'b0;
    assign data[2833] = ~16'b0;
    assign data[2834] = ~16'b0;
    assign data[2835] = ~16'b0;
    assign data[2836] = ~16'b0;
    assign data[2837] = ~16'b0;
    assign data[2838] = ~16'b0;
    assign data[2839] = ~16'b0;
    assign data[2840] = 16'b0;
    assign data[2841] = 16'b0;
    assign data[2842] = ~16'b0;
    assign data[2843] = ~16'b0;
    assign data[2844] = ~16'b0;
    assign data[2845] = ~16'b0;
    assign data[2846] = ~16'b0;
    assign data[2847] = ~16'b0;
    assign data[2848] = ~16'b0;
    assign data[2849] = ~16'b0;
    assign data[2850] = 16'b0;
    assign data[2851] = 16'b0;
    assign data[2852] = ~16'b0;
    assign data[2853] = ~16'b0;
    assign data[2854] = ~16'b0;
    assign data[2855] = ~16'b0;
    assign data[2856] = ~16'b0;
    assign data[2857] = ~16'b0;
    assign data[2858] = ~16'b0;
    assign data[2859] = ~16'b0;
    assign data[2860] = 16'b0;
    assign data[2861] = 16'b0;
    assign data[2862] = ~16'b0;
    assign data[2863] = ~16'b0;
    assign data[2864] = ~16'b0;
    assign data[2865] = ~16'b0;
    assign data[2866] = ~16'b0;
    assign data[2867] = ~16'b0;
    assign data[2868] = ~16'b0;
    assign data[2869] = ~16'b0;
    assign data[2870] = 16'b0;
    assign data[2871] = 16'b0;
    assign data[2872] = ~16'b0;
    assign data[2873] = ~16'b0;
    assign data[2874] = ~16'b0;
    assign data[2875] = ~16'b0;
    assign data[2876] = ~16'b0;
    assign data[2877] = ~16'b0;
    assign data[2878] = ~16'b0;
    assign data[2879] = ~16'b0;
    assign data[2880] = 16'b0;
    assign data[2881] = 16'b0;
    assign data[2882] = ~16'b0;
    assign data[2883] = ~16'b0;
    assign data[2884] = ~16'b0;
    assign data[2885] = ~16'b0;
    assign data[2886] = ~16'b0;
    assign data[2887] = ~16'b0;
    assign data[2888] = ~16'b0;
    assign data[2889] = ~16'b0;
    assign data[2890] = 16'b0;
    assign data[2891] = 16'b0;
    assign data[2892] = ~16'b0;
    assign data[2893] = ~16'b0;
    assign data[2894] = ~16'b0;
    assign data[2895] = ~16'b0;
    assign data[2896] = ~16'b0;
    assign data[2897] = ~16'b0;
    assign data[2898] = ~16'b0;
    assign data[2899] = ~16'b0;
    assign data[2900] = 16'b0;
    assign data[2901] = 16'b0;
    assign data[2902] = ~16'b0;
    assign data[2903] = ~16'b0;
    assign data[2904] = ~16'b0;
    assign data[2905] = ~16'b0;
    assign data[2906] = ~16'b0;
    assign data[2907] = ~16'b0;
    assign data[2908] = ~16'b0;
    assign data[2909] = ~16'b0;
    assign data[2910] = 16'b0;
    assign data[2911] = 16'b0;
    assign data[2912] = ~16'b0;
    assign data[2913] = ~16'b0;
    assign data[2914] = ~16'b0;
    assign data[2915] = ~16'b0;
    assign data[2916] = ~16'b0;
    assign data[2917] = ~16'b0;
    assign data[2918] = ~16'b0;
    assign data[2919] = ~16'b0;
    assign data[2920] = 16'b0;
    assign data[2921] = 16'b0;
    assign data[2922] = ~16'b0;
    assign data[2923] = ~16'b0;
    assign data[2924] = ~16'b0;
    assign data[2925] = ~16'b0;
    assign data[2926] = ~16'b0;
    assign data[2927] = ~16'b0;
    assign data[2928] = ~16'b0;
    assign data[2929] = ~16'b0;
    assign data[2930] = 16'b0;
    assign data[2931] = 16'b0;
    assign data[2932] = ~16'b0;
    assign data[2933] = ~16'b0;
    assign data[2934] = ~16'b0;
    assign data[2935] = ~16'b0;
    assign data[2936] = ~16'b0;
    assign data[2937] = ~16'b0;
    assign data[2938] = ~16'b0;
    assign data[2939] = ~16'b0;
    assign data[2940] = 16'b0;
    assign data[2941] = 16'b0;
    assign data[2942] = ~16'b0;
    assign data[2943] = ~16'b0;
    assign data[2944] = ~16'b0;
    assign data[2945] = ~16'b0;
    assign data[2946] = ~16'b0;
    assign data[2947] = ~16'b0;
    assign data[2948] = ~16'b0;
    assign data[2949] = ~16'b0;
    assign data[2950] = 16'b0;
    assign data[2951] = 16'b0;
    assign data[2952] = ~16'b0;
    assign data[2953] = ~16'b0;
    assign data[2954] = ~16'b0;
    assign data[2955] = ~16'b0;
    assign data[2956] = ~16'b0;
    assign data[2957] = ~16'b0;
    assign data[2958] = ~16'b0;
    assign data[2959] = ~16'b0;
    assign data[2960] = 16'b0;
    assign data[2961] = 16'b0;
    assign data[2962] = ~16'b0;
    assign data[2963] = ~16'b0;
    assign data[2964] = ~16'b0;
    assign data[2965] = ~16'b0;
    assign data[2966] = ~16'b0;
    assign data[2967] = ~16'b0;
    assign data[2968] = ~16'b0;
    assign data[2969] = ~16'b0;
    assign data[2970] = 16'b0;
    assign data[2971] = 16'b0;
    assign data[2972] = ~16'b0;
    assign data[2973] = ~16'b0;
    assign data[2974] = ~16'b0;
    assign data[2975] = ~16'b0;
    assign data[2976] = ~16'b0;
    assign data[2977] = ~16'b0;
    assign data[2978] = ~16'b0;
    assign data[2979] = ~16'b0;
    assign data[2980] = 16'b0;
    assign data[2981] = 16'b0;
    assign data[2982] = ~16'b0;
    assign data[2983] = ~16'b0;
    assign data[2984] = ~16'b0;
    assign data[2985] = ~16'b0;
    assign data[2986] = ~16'b0;
    assign data[2987] = ~16'b0;
    assign data[2988] = ~16'b0;
    assign data[2989] = ~16'b0;
    assign data[2990] = 16'b0;
    assign data[2991] = 16'b0;
    assign data[2992] = ~16'b0;
    assign data[2993] = ~16'b0;
    assign data[2994] = ~16'b0;
    assign data[2995] = ~16'b0;
    assign data[2996] = ~16'b0;
    assign data[2997] = ~16'b0;
    assign data[2998] = ~16'b0;
    assign data[2999] = ~16'b0;
    assign data[3000] = 16'b0;
    assign data[3001] = 16'b0;
    assign data[3002] = ~16'b0;
    assign data[3003] = ~16'b0;
    assign data[3004] = ~16'b0;
    assign data[3005] = ~16'b0;
    assign data[3006] = ~16'b0;
    assign data[3007] = ~16'b0;
    assign data[3008] = ~16'b0;
    assign data[3009] = ~16'b0;
    assign data[3010] = 16'b0;
    assign data[3011] = 16'b0;
    assign data[3012] = 16'b0;
    assign data[3013] = 16'b0;
    assign data[3014] = 16'b0;
    assign data[3015] = 16'b0;
    assign data[3016] = 16'b0;
    assign data[3017] = 16'b0;
    assign data[3018] = 16'b0;
    assign data[3019] = 16'b0;
    assign data[3020] = 16'b0;
    assign data[3021] = 16'b0;
    assign data[3022] = 16'b0;
    assign data[3023] = 16'b0;
    assign data[3024] = 16'b0;
    assign data[3025] = 16'b0;
    assign data[3026] = 16'b0;
    assign data[3027] = 16'b0;
    assign data[3028] = 16'b0;
    assign data[3029] = 16'b0;
    assign data[3030] = ~16'b0;
    assign data[3031] = ~16'b0;
    assign data[3032] = ~16'b0;
    assign data[3033] = ~16'b0;
    assign data[3034] = ~16'b0;
    assign data[3035] = ~16'b0;
    assign data[3036] = ~16'b0;
    assign data[3037] = ~16'b0;
    assign data[3038] = ~16'b0;
    assign data[3039] = ~16'b0;
    assign data[3040] = ~16'b0;
    assign data[3041] = ~16'b0;
    assign data[3042] = ~16'b0;
    assign data[3043] = ~16'b0;
    assign data[3044] = ~16'b0;
    assign data[3045] = ~16'b0;
    assign data[3046] = ~16'b0;
    assign data[3047] = ~16'b0;
    assign data[3048] = ~16'b0;
    assign data[3049] = ~16'b0;
    assign data[3050] = ~16'b0;
    assign data[3051] = ~16'b0;
    assign data[3052] = ~16'b0;
    assign data[3053] = ~16'b0;
    assign data[3054] = ~16'b0;
    assign data[3055] = ~16'b0;
    assign data[3056] = ~16'b0;
    assign data[3057] = ~16'b0;
    assign data[3058] = ~16'b0;
    assign data[3059] = ~16'b0;
    assign data[3060] = ~16'b0;
    assign data[3061] = ~16'b0;
    assign data[3062] = ~16'b0;
    assign data[3063] = ~16'b0;
    assign data[3064] = ~16'b0;
    assign data[3065] = ~16'b0;
    assign data[3066] = ~16'b0;
    assign data[3067] = ~16'b0;
    assign data[3068] = ~16'b0;
    assign data[3069] = ~16'b0;
    assign data[3070] = ~16'b0;
    assign data[3071] = ~16'b0;
    assign data[3072] = ~16'b0;
    assign data[3073] = ~16'b0;
    assign data[3074] = ~16'b0;
    assign data[3075] = ~16'b0;
    assign data[3076] = ~16'b0;
    assign data[3077] = ~16'b0;
    assign data[3078] = ~16'b0;
    assign data[3079] = ~16'b0;
    assign data[3080] = ~16'b0;
    assign data[3081] = ~16'b0;
    assign data[3082] = ~16'b0;
    assign data[3083] = ~16'b0;
    assign data[3084] = ~16'b0;
    assign data[3085] = ~16'b0;
    assign data[3086] = ~16'b0;
    assign data[3087] = ~16'b0;
    assign data[3088] = ~16'b0;
    assign data[3089] = ~16'b0;
    assign data[3090] = ~16'b0;
    assign data[3091] = ~16'b0;
    assign data[3092] = ~16'b0;
    assign data[3093] = ~16'b0;
    assign data[3094] = ~16'b0;
    assign data[3095] = ~16'b0;
    assign data[3096] = ~16'b0;
    assign data[3097] = ~16'b0;
    assign data[3098] = ~16'b0;
    assign data[3099] = ~16'b0;
    assign data[3100] = ~16'b0;
    assign data[3101] = ~16'b0;
    assign data[3102] = ~16'b0;
    assign data[3103] = ~16'b0;
    assign data[3104] = ~16'b0;
    assign data[3105] = ~16'b0;
    assign data[3106] = ~16'b0;
    assign data[3107] = ~16'b0;
    assign data[3108] = ~16'b0;
    assign data[3109] = ~16'b0;
    assign data[3110] = ~16'b0;
    assign data[3111] = ~16'b0;
    assign data[3112] = ~16'b0;
    assign data[3113] = ~16'b0;
    assign data[3114] = ~16'b0;
    assign data[3115] = ~16'b0;
    assign data[3116] = ~16'b0;
    assign data[3117] = ~16'b0;
    assign data[3118] = ~16'b0;
    assign data[3119] = ~16'b0;
    assign data[3120] = ~16'b0;
    assign data[3121] = ~16'b0;
    assign data[3122] = ~16'b0;
    assign data[3123] = ~16'b0;
    assign data[3124] = ~16'b0;
    assign data[3125] = ~16'b0;
    assign data[3126] = ~16'b0;
    assign data[3127] = ~16'b0;
    assign data[3128] = ~16'b0;
    assign data[3129] = ~16'b0;
    assign data[3130] = ~16'b0;
    assign data[3131] = ~16'b0;
    assign data[3132] = ~16'b0;
    assign data[3133] = ~16'b0;
    assign data[3134] = ~16'b0;
    assign data[3135] = ~16'b0;
    assign data[3136] = ~16'b0;
    assign data[3137] = ~16'b0;
    assign data[3138] = ~16'b0;
    assign data[3139] = ~16'b0;
    assign data[3140] = ~16'b0;
    assign data[3141] = ~16'b0;
    assign data[3142] = ~16'b0;
    assign data[3143] = ~16'b0;
    assign data[3144] = ~16'b0;
    assign data[3145] = ~16'b0;
    assign data[3146] = ~16'b0;
    assign data[3147] = ~16'b0;
    assign data[3148] = ~16'b0;
    assign data[3149] = ~16'b0;
    assign data[3150] = ~16'b0;
    assign data[3151] = ~16'b0;
    assign data[3152] = ~16'b0;
    assign data[3153] = ~16'b0;
    assign data[3154] = ~16'b0;
    assign data[3155] = ~16'b0;
    assign data[3156] = ~16'b0;
    assign data[3157] = ~16'b0;
    assign data[3158] = ~16'b0;
    assign data[3159] = ~16'b0;
    assign data[3160] = ~16'b0;
    assign data[3161] = ~16'b0;
    assign data[3162] = ~16'b0;
    assign data[3163] = ~16'b0;
    assign data[3164] = ~16'b0;
    assign data[3165] = ~16'b0;
    assign data[3166] = ~16'b0;
    assign data[3167] = ~16'b0;
    assign data[3168] = ~16'b0;
    assign data[3169] = ~16'b0;
    assign data[3170] = ~16'b0;
    assign data[3171] = ~16'b0;
    assign data[3172] = ~16'b0;
    assign data[3173] = ~16'b0;
    assign data[3174] = ~16'b0;
    assign data[3175] = ~16'b0;
    assign data[3176] = ~16'b0;
    assign data[3177] = ~16'b0;
    assign data[3178] = ~16'b0;
    assign data[3179] = ~16'b0;
    assign data[3180] = ~16'b0;
    assign data[3181] = ~16'b0;
    assign data[3182] = ~16'b0;
    assign data[3183] = ~16'b0;
    assign data[3184] = ~16'b0;
    assign data[3185] = ~16'b0;
    assign data[3186] = ~16'b0;
    assign data[3187] = ~16'b0;
    assign data[3188] = ~16'b0;
    assign data[3189] = ~16'b0;
    assign data[3190] = ~16'b0;
    assign data[3191] = ~16'b0;
    assign data[3192] = ~16'b0;
    assign data[3193] = ~16'b0;
    assign data[3194] = ~16'b0;
    assign data[3195] = ~16'b0;
    assign data[3196] = ~16'b0;
    assign data[3197] = ~16'b0;
    assign data[3198] = ~16'b0;
    assign data[3199] = ~16'b0;
    assign data[3200] = ~16'b0;
    assign data[3201] = ~16'b0;
    assign data[3202] = ~16'b0;
    assign data[3203] = ~16'b0;
    assign data[3204] = ~16'b0;
    assign data[3205] = ~16'b0;
    assign data[3206] = ~16'b0;
    assign data[3207] = ~16'b0;
    assign data[3208] = ~16'b0;
    assign data[3209] = ~16'b0;
    assign data[3210] = ~16'b0;
    assign data[3211] = ~16'b0;
    assign data[3212] = ~16'b0;
    assign data[3213] = ~16'b0;
    assign data[3214] = ~16'b0;
    assign data[3215] = ~16'b0;
    assign data[3216] = ~16'b0;
    assign data[3217] = ~16'b0;
    assign data[3218] = ~16'b0;
    assign data[3219] = ~16'b0;
    assign data[3220] = ~16'b0;
    assign data[3221] = ~16'b0;
    assign data[3222] = ~16'b0;
    assign data[3223] = ~16'b0;
    assign data[3224] = ~16'b0;
    assign data[3225] = ~16'b0;
    assign data[3226] = ~16'b0;
    assign data[3227] = ~16'b0;
    assign data[3228] = ~16'b0;
    assign data[3229] = ~16'b0;
    assign data[3230] = ~16'b0;
    assign data[3231] = ~16'b0;
    assign data[3232] = ~16'b0;
    assign data[3233] = ~16'b0;
    assign data[3234] = ~16'b0;
    assign data[3235] = ~16'b0;
    assign data[3236] = ~16'b0;
    assign data[3237] = ~16'b0;
    assign data[3238] = ~16'b0;
    assign data[3239] = ~16'b0;
    assign data[3240] = ~16'b0;
    assign data[3241] = ~16'b0;
    assign data[3242] = ~16'b0;
    assign data[3243] = ~16'b0;
    assign data[3244] = ~16'b0;
    assign data[3245] = ~16'b0;
    assign data[3246] = ~16'b0;
    assign data[3247] = ~16'b0;
    assign data[3248] = ~16'b0;
    assign data[3249] = ~16'b0;
    assign data[3250] = ~16'b0;
    assign data[3251] = ~16'b0;
    assign data[3252] = ~16'b0;
    assign data[3253] = ~16'b0;
    assign data[3254] = ~16'b0;
    assign data[3255] = ~16'b0;
    assign data[3256] = ~16'b0;
    assign data[3257] = ~16'b0;
    assign data[3258] = ~16'b0;
    assign data[3259] = ~16'b0;
    assign data[3260] = ~16'b0;
    assign data[3261] = ~16'b0;
    assign data[3262] = ~16'b0;
    assign data[3263] = ~16'b0;
    assign data[3264] = ~16'b0;
    assign data[3265] = ~16'b0;
    assign data[3266] = ~16'b0;
    assign data[3267] = ~16'b0;
    assign data[3268] = ~16'b0;
    assign data[3269] = ~16'b0;
    assign data[3270] = 16'b0;
    assign data[3271] = 16'b0;
    assign data[3272] = 16'b0;
    assign data[3273] = 16'b0;
    assign data[3274] = 16'b0;
    assign data[3275] = 16'b0;
    assign data[3276] = 16'b0;
    assign data[3277] = 16'b0;
    assign data[3278] = 16'b0;
    assign data[3279] = 16'b0;
    assign data[3280] = 16'b0;
    assign data[3281] = 16'b0;
    assign data[3282] = 16'b0;
    assign data[3283] = 16'b0;
    assign data[3284] = 16'b0;
    assign data[3285] = 16'b0;
    assign data[3286] = 16'b0;
    assign data[3287] = 16'b0;
    assign data[3288] = 16'b0;
    assign data[3289] = 16'b0;
    assign data[3290] = 16'b0;
    assign data[3291] = 16'b0;
    assign data[3292] = ~16'b0;
    assign data[3293] = ~16'b0;
    assign data[3294] = ~16'b0;
    assign data[3295] = ~16'b0;
    assign data[3296] = ~16'b0;
    assign data[3297] = ~16'b0;
    assign data[3298] = ~16'b0;
    assign data[3299] = ~16'b0;
    assign data[3300] = 16'b0;
    assign data[3301] = 16'b0;
    assign data[3302] = ~16'b0;
    assign data[3303] = ~16'b0;
    assign data[3304] = ~16'b0;
    assign data[3305] = ~16'b0;
    assign data[3306] = ~16'b0;
    assign data[3307] = ~16'b0;
    assign data[3308] = ~16'b0;
    assign data[3309] = ~16'b0;
    assign data[3310] = 16'b0;
    assign data[3311] = 16'b0;
    assign data[3312] = ~16'b0;
    assign data[3313] = ~16'b0;
    assign data[3314] = ~16'b0;
    assign data[3315] = ~16'b0;
    assign data[3316] = ~16'b0;
    assign data[3317] = ~16'b0;
    assign data[3318] = ~16'b0;
    assign data[3319] = ~16'b0;
    assign data[3320] = 16'b0;
    assign data[3321] = 16'b0;
    assign data[3322] = ~16'b0;
    assign data[3323] = ~16'b0;
    assign data[3324] = ~16'b0;
    assign data[3325] = ~16'b0;
    assign data[3326] = ~16'b0;
    assign data[3327] = ~16'b0;
    assign data[3328] = ~16'b0;
    assign data[3329] = ~16'b0;
    assign data[3330] = 16'b0;
    assign data[3331] = 16'b0;
    assign data[3332] = ~16'b0;
    assign data[3333] = ~16'b0;
    assign data[3334] = ~16'b0;
    assign data[3335] = ~16'b0;
    assign data[3336] = ~16'b0;
    assign data[3337] = ~16'b0;
    assign data[3338] = ~16'b0;
    assign data[3339] = ~16'b0;
    assign data[3340] = 16'b0;
    assign data[3341] = 16'b0;
    assign data[3342] = ~16'b0;
    assign data[3343] = ~16'b0;
    assign data[3344] = ~16'b0;
    assign data[3345] = ~16'b0;
    assign data[3346] = ~16'b0;
    assign data[3347] = ~16'b0;
    assign data[3348] = ~16'b0;
    assign data[3349] = ~16'b0;
    assign data[3350] = 16'b0;
    assign data[3351] = 16'b0;
    assign data[3352] = ~16'b0;
    assign data[3353] = ~16'b0;
    assign data[3354] = ~16'b0;
    assign data[3355] = ~16'b0;
    assign data[3356] = ~16'b0;
    assign data[3357] = ~16'b0;
    assign data[3358] = ~16'b0;
    assign data[3359] = ~16'b0;
    assign data[3360] = 16'b0;
    assign data[3361] = 16'b0;
    assign data[3362] = ~16'b0;
    assign data[3363] = ~16'b0;
    assign data[3364] = ~16'b0;
    assign data[3365] = ~16'b0;
    assign data[3366] = ~16'b0;
    assign data[3367] = ~16'b0;
    assign data[3368] = ~16'b0;
    assign data[3369] = ~16'b0;
    assign data[3370] = 16'b0;
    assign data[3371] = 16'b0;
    assign data[3372] = ~16'b0;
    assign data[3373] = ~16'b0;
    assign data[3374] = ~16'b0;
    assign data[3375] = ~16'b0;
    assign data[3376] = ~16'b0;
    assign data[3377] = ~16'b0;
    assign data[3378] = ~16'b0;
    assign data[3379] = ~16'b0;
    assign data[3380] = 16'b0;
    assign data[3381] = 16'b0;
    assign data[3382] = ~16'b0;
    assign data[3383] = ~16'b0;
    assign data[3384] = ~16'b0;
    assign data[3385] = ~16'b0;
    assign data[3386] = ~16'b0;
    assign data[3387] = ~16'b0;
    assign data[3388] = ~16'b0;
    assign data[3389] = ~16'b0;
    assign data[3390] = 16'b0;
    assign data[3391] = 16'b0;
    assign data[3392] = ~16'b0;
    assign data[3393] = ~16'b0;
    assign data[3394] = ~16'b0;
    assign data[3395] = ~16'b0;
    assign data[3396] = ~16'b0;
    assign data[3397] = ~16'b0;
    assign data[3398] = ~16'b0;
    assign data[3399] = ~16'b0;
    assign data[3400] = 16'b0;
    assign data[3401] = 16'b0;
    assign data[3402] = ~16'b0;
    assign data[3403] = ~16'b0;
    assign data[3404] = ~16'b0;
    assign data[3405] = ~16'b0;
    assign data[3406] = ~16'b0;
    assign data[3407] = ~16'b0;
    assign data[3408] = ~16'b0;
    assign data[3409] = ~16'b0;
    assign data[3410] = 16'b0;
    assign data[3411] = 16'b0;
    assign data[3412] = ~16'b0;
    assign data[3413] = ~16'b0;
    assign data[3414] = ~16'b0;
    assign data[3415] = ~16'b0;
    assign data[3416] = ~16'b0;
    assign data[3417] = ~16'b0;
    assign data[3418] = ~16'b0;
    assign data[3419] = ~16'b0;
    assign data[3420] = 16'b0;
    assign data[3421] = 16'b0;
    assign data[3422] = ~16'b0;
    assign data[3423] = ~16'b0;
    assign data[3424] = ~16'b0;
    assign data[3425] = ~16'b0;
    assign data[3426] = ~16'b0;
    assign data[3427] = ~16'b0;
    assign data[3428] = ~16'b0;
    assign data[3429] = ~16'b0;
    assign data[3430] = 16'b0;
    assign data[3431] = 16'b0;
    assign data[3432] = ~16'b0;
    assign data[3433] = ~16'b0;
    assign data[3434] = ~16'b0;
    assign data[3435] = ~16'b0;
    assign data[3436] = ~16'b0;
    assign data[3437] = ~16'b0;
    assign data[3438] = ~16'b0;
    assign data[3439] = ~16'b0;
    assign data[3440] = 16'b0;
    assign data[3441] = 16'b0;
    assign data[3442] = ~16'b0;
    assign data[3443] = ~16'b0;
    assign data[3444] = ~16'b0;
    assign data[3445] = ~16'b0;
    assign data[3446] = ~16'b0;
    assign data[3447] = ~16'b0;
    assign data[3448] = ~16'b0;
    assign data[3449] = ~16'b0;
    assign data[3450] = 16'b0;
    assign data[3451] = 16'b0;
    assign data[3452] = ~16'b0;
    assign data[3453] = ~16'b0;
    assign data[3454] = ~16'b0;
    assign data[3455] = ~16'b0;
    assign data[3456] = ~16'b0;
    assign data[3457] = ~16'b0;
    assign data[3458] = ~16'b0;
    assign data[3459] = ~16'b0;
    assign data[3460] = 16'b0;
    assign data[3461] = 16'b0;
    assign data[3462] = ~16'b0;
    assign data[3463] = ~16'b0;
    assign data[3464] = ~16'b0;
    assign data[3465] = ~16'b0;
    assign data[3466] = ~16'b0;
    assign data[3467] = ~16'b0;
    assign data[3468] = ~16'b0;
    assign data[3469] = ~16'b0;
    assign data[3470] = 16'b0;
    assign data[3471] = 16'b0;
    assign data[3472] = ~16'b0;
    assign data[3473] = ~16'b0;
    assign data[3474] = ~16'b0;
    assign data[3475] = ~16'b0;
    assign data[3476] = ~16'b0;
    assign data[3477] = ~16'b0;
    assign data[3478] = ~16'b0;
    assign data[3479] = ~16'b0;
    assign data[3480] = 16'b0;
    assign data[3481] = 16'b0;
    assign data[3482] = ~16'b0;
    assign data[3483] = ~16'b0;
    assign data[3484] = ~16'b0;
    assign data[3485] = ~16'b0;
    assign data[3486] = ~16'b0;
    assign data[3487] = ~16'b0;
    assign data[3488] = ~16'b0;
    assign data[3489] = ~16'b0;
    assign data[3490] = 16'b0;
    assign data[3491] = 16'b0;
    assign data[3492] = ~16'b0;
    assign data[3493] = ~16'b0;
    assign data[3494] = ~16'b0;
    assign data[3495] = ~16'b0;
    assign data[3496] = ~16'b0;
    assign data[3497] = ~16'b0;
    assign data[3498] = ~16'b0;
    assign data[3499] = ~16'b0;
    assign data[3500] = 16'b0;
    assign data[3501] = 16'b0;
    assign data[3502] = ~16'b0;
    assign data[3503] = ~16'b0;
    assign data[3504] = ~16'b0;
    assign data[3505] = ~16'b0;
    assign data[3506] = ~16'b0;
    assign data[3507] = ~16'b0;
    assign data[3508] = ~16'b0;
    assign data[3509] = ~16'b0;
    assign data[3510] = 16'b0;
    assign data[3511] = 16'b0;
    assign data[3512] = ~16'b0;
    assign data[3513] = ~16'b0;
    assign data[3514] = ~16'b0;
    assign data[3515] = ~16'b0;
    assign data[3516] = ~16'b0;
    assign data[3517] = ~16'b0;
    assign data[3518] = ~16'b0;
    assign data[3519] = ~16'b0;
    assign data[3520] = 16'b0;
    assign data[3521] = 16'b0;
    assign data[3522] = ~16'b0;
    assign data[3523] = ~16'b0;
    assign data[3524] = ~16'b0;
    assign data[3525] = ~16'b0;
    assign data[3526] = ~16'b0;
    assign data[3527] = ~16'b0;
    assign data[3528] = ~16'b0;
    assign data[3529] = ~16'b0;
    assign data[3530] = 16'b0;
    assign data[3531] = 16'b0;
    assign data[3532] = ~16'b0;
    assign data[3533] = ~16'b0;
    assign data[3534] = ~16'b0;
    assign data[3535] = ~16'b0;
    assign data[3536] = ~16'b0;
    assign data[3537] = ~16'b0;
    assign data[3538] = ~16'b0;
    assign data[3539] = ~16'b0;
    assign data[3540] = 16'b0;
    assign data[3541] = 16'b0;
    assign data[3542] = ~16'b0;
    assign data[3543] = ~16'b0;
    assign data[3544] = ~16'b0;
    assign data[3545] = ~16'b0;
    assign data[3546] = ~16'b0;
    assign data[3547] = ~16'b0;
    assign data[3548] = ~16'b0;
    assign data[3549] = ~16'b0;
    assign data[3550] = 16'b0;
    assign data[3551] = 16'b0;
    assign data[3552] = ~16'b0;
    assign data[3553] = ~16'b0;
    assign data[3554] = ~16'b0;
    assign data[3555] = ~16'b0;
    assign data[3556] = ~16'b0;
    assign data[3557] = ~16'b0;
    assign data[3558] = ~16'b0;
    assign data[3559] = ~16'b0;
    assign data[3560] = 16'b0;
    assign data[3561] = 16'b0;
    assign data[3562] = ~16'b0;
    assign data[3563] = ~16'b0;
    assign data[3564] = ~16'b0;
    assign data[3565] = ~16'b0;
    assign data[3566] = ~16'b0;
    assign data[3567] = ~16'b0;
    assign data[3568] = ~16'b0;
    assign data[3569] = ~16'b0;
    assign data[3570] = 16'b0;
    assign data[3571] = 16'b0;
    assign data[3572] = ~16'b0;
    assign data[3573] = ~16'b0;
    assign data[3574] = ~16'b0;
    assign data[3575] = ~16'b0;
    assign data[3576] = ~16'b0;
    assign data[3577] = ~16'b0;
    assign data[3578] = ~16'b0;
    assign data[3579] = ~16'b0;
    assign data[3580] = 16'b0;
    assign data[3581] = 16'b0;
    assign data[3582] = ~16'b0;
    assign data[3583] = ~16'b0;
    assign data[3584] = ~16'b0;
    assign data[3585] = ~16'b0;
    assign data[3586] = ~16'b0;
    assign data[3587] = ~16'b0;
    assign data[3588] = ~16'b0;
    assign data[3589] = ~16'b0;
    assign data[3590] = 16'b0;
    assign data[3591] = 16'b0;
    assign data[3592] = ~16'b0;
    assign data[3593] = ~16'b0;
    assign data[3594] = ~16'b0;
    assign data[3595] = ~16'b0;
    assign data[3596] = ~16'b0;
    assign data[3597] = ~16'b0;
    assign data[3598] = ~16'b0;
    assign data[3599] = ~16'b0;
    assign data[3600] = 16'b0;
    assign data[3601] = 16'b0;
    assign data[3602] = ~16'b0;
    assign data[3603] = ~16'b0;
    assign data[3604] = ~16'b0;
    assign data[3605] = ~16'b0;
    assign data[3606] = ~16'b0;
    assign data[3607] = ~16'b0;
    assign data[3608] = ~16'b0;
    assign data[3609] = ~16'b0;
    assign data[3610] = 16'b0;
    assign data[3611] = 16'b0;
    assign data[3612] = 16'b0;
    assign data[3613] = 16'b0;
    assign data[3614] = 16'b0;
    assign data[3615] = 16'b0;
    assign data[3616] = 16'b0;
    assign data[3617] = 16'b0;
    assign data[3618] = 16'b0;
    assign data[3619] = 16'b0;
    assign data[3620] = 16'b0;
    assign data[3621] = 16'b0;
    assign data[3622] = 16'b0;
    assign data[3623] = 16'b0;
    assign data[3624] = 16'b0;
    assign data[3625] = 16'b0;
    assign data[3626] = 16'b0;
    assign data[3627] = 16'b0;
    assign data[3628] = 16'b0;
    assign data[3629] = 16'b0;
    assign data[3630] = ~16'b0;
    assign data[3631] = ~16'b0;
    assign data[3632] = ~16'b0;
    assign data[3633] = ~16'b0;
    assign data[3634] = ~16'b0;
    assign data[3635] = ~16'b0;
    assign data[3636] = ~16'b0;
    assign data[3637] = ~16'b0;
    assign data[3638] = ~16'b0;
    assign data[3639] = ~16'b0;
    assign data[3640] = ~16'b0;
    assign data[3641] = ~16'b0;
    assign data[3642] = ~16'b0;
    assign data[3643] = ~16'b0;
    assign data[3644] = ~16'b0;
    assign data[3645] = ~16'b0;
    assign data[3646] = ~16'b0;
    assign data[3647] = ~16'b0;
    assign data[3648] = ~16'b0;
    assign data[3649] = ~16'b0;
    assign data[3650] = ~16'b0;
    assign data[3651] = ~16'b0;
    assign data[3652] = ~16'b0;
    assign data[3653] = ~16'b0;
    assign data[3654] = ~16'b0;
    assign data[3655] = ~16'b0;
    assign data[3656] = ~16'b0;
    assign data[3657] = ~16'b0;
    assign data[3658] = ~16'b0;
    assign data[3659] = ~16'b0;
    assign data[3660] = ~16'b0;
    assign data[3661] = ~16'b0;
    assign data[3662] = ~16'b0;
    assign data[3663] = ~16'b0;
    assign data[3664] = ~16'b0;
    assign data[3665] = ~16'b0;
    assign data[3666] = ~16'b0;
    assign data[3667] = ~16'b0;
    assign data[3668] = ~16'b0;
    assign data[3669] = ~16'b0;
    assign data[3670] = ~16'b0;
    assign data[3671] = ~16'b0;
    assign data[3672] = ~16'b0;
    assign data[3673] = ~16'b0;
    assign data[3674] = ~16'b0;
    assign data[3675] = ~16'b0;
    assign data[3676] = ~16'b0;
    assign data[3677] = ~16'b0;
    assign data[3678] = ~16'b0;
    assign data[3679] = ~16'b0;
    assign data[3680] = ~16'b0;
    assign data[3681] = ~16'b0;
    assign data[3682] = ~16'b0;
    assign data[3683] = ~16'b0;
    assign data[3684] = ~16'b0;
    assign data[3685] = ~16'b0;
    assign data[3686] = ~16'b0;
    assign data[3687] = ~16'b0;
    assign data[3688] = ~16'b0;
    assign data[3689] = ~16'b0;
    assign data[3690] = ~16'b0;
    assign data[3691] = ~16'b0;
    assign data[3692] = ~16'b0;
    assign data[3693] = ~16'b0;
    assign data[3694] = ~16'b0;
    assign data[3695] = ~16'b0;
    assign data[3696] = ~16'b0;
    assign data[3697] = ~16'b0;
    assign data[3698] = ~16'b0;
    assign data[3699] = ~16'b0;
    assign data[3700] = ~16'b0;
    assign data[3701] = ~16'b0;
    assign data[3702] = ~16'b0;
    assign data[3703] = ~16'b0;
    assign data[3704] = ~16'b0;
    assign data[3705] = ~16'b0;
    assign data[3706] = ~16'b0;
    assign data[3707] = ~16'b0;
    assign data[3708] = ~16'b0;
    assign data[3709] = ~16'b0;
    assign data[3710] = ~16'b0;
    assign data[3711] = ~16'b0;
    assign data[3712] = ~16'b0;
    assign data[3713] = ~16'b0;
    assign data[3714] = ~16'b0;
    assign data[3715] = ~16'b0;
    assign data[3716] = ~16'b0;
    assign data[3717] = ~16'b0;
    assign data[3718] = ~16'b0;
    assign data[3719] = ~16'b0;
    assign data[3720] = ~16'b0;
    assign data[3721] = ~16'b0;
    assign data[3722] = ~16'b0;
    assign data[3723] = ~16'b0;
    assign data[3724] = ~16'b0;
    assign data[3725] = ~16'b0;
    assign data[3726] = ~16'b0;
    assign data[3727] = ~16'b0;
    assign data[3728] = ~16'b0;
    assign data[3729] = ~16'b0;
    assign data[3730] = ~16'b0;
    assign data[3731] = ~16'b0;
    assign data[3732] = ~16'b0;
    assign data[3733] = ~16'b0;
    assign data[3734] = ~16'b0;
    assign data[3735] = ~16'b0;
    assign data[3736] = ~16'b0;
    assign data[3737] = ~16'b0;
    assign data[3738] = ~16'b0;
    assign data[3739] = ~16'b0;
    assign data[3740] = ~16'b0;
    assign data[3741] = ~16'b0;
    assign data[3742] = ~16'b0;
    assign data[3743] = ~16'b0;
    assign data[3744] = ~16'b0;
    assign data[3745] = ~16'b0;
    assign data[3746] = ~16'b0;
    assign data[3747] = ~16'b0;
    assign data[3748] = ~16'b0;
    assign data[3749] = ~16'b0;
    assign data[3750] = ~16'b0;
    assign data[3751] = ~16'b0;
    assign data[3752] = ~16'b0;
    assign data[3753] = ~16'b0;
    assign data[3754] = ~16'b0;
    assign data[3755] = ~16'b0;
    assign data[3756] = ~16'b0;
    assign data[3757] = ~16'b0;
    assign data[3758] = ~16'b0;
    assign data[3759] = ~16'b0;
    assign data[3760] = ~16'b0;
    assign data[3761] = ~16'b0;
    assign data[3762] = ~16'b0;
    assign data[3763] = ~16'b0;
    assign data[3764] = ~16'b0;
    assign data[3765] = ~16'b0;
    assign data[3766] = ~16'b0;
    assign data[3767] = ~16'b0;
    assign data[3768] = ~16'b0;
    assign data[3769] = ~16'b0;
    assign data[3770] = ~16'b0;
    assign data[3771] = ~16'b0;
    assign data[3772] = ~16'b0;
    assign data[3773] = ~16'b0;
    assign data[3774] = ~16'b0;
    assign data[3775] = ~16'b0;
    assign data[3776] = ~16'b0;
    assign data[3777] = ~16'b0;
    assign data[3778] = ~16'b0;
    assign data[3779] = ~16'b0;
    assign data[3780] = ~16'b0;
    assign data[3781] = ~16'b0;
    assign data[3782] = ~16'b0;
    assign data[3783] = ~16'b0;
    assign data[3784] = ~16'b0;
    assign data[3785] = ~16'b0;
    assign data[3786] = ~16'b0;
    assign data[3787] = ~16'b0;
    assign data[3788] = ~16'b0;
    assign data[3789] = ~16'b0;
    assign data[3790] = 16'b0;
    assign data[3791] = 16'b0;
    assign data[3792] = 16'b0;
    assign data[3793] = 16'b0;
    assign data[3794] = 16'b0;
    assign data[3795] = 16'b0;
    assign data[3796] = 16'b0;
    assign data[3797] = 16'b0;
    assign data[3798] = 16'b0;
    assign data[3799] = 16'b0;
    assign data[3800] = 16'b0;
    assign data[3801] = 16'b0;
    assign data[3802] = 16'b0;
    assign data[3803] = 16'b0;
    assign data[3804] = 16'b0;
    assign data[3805] = 16'b0;
    assign data[3806] = 16'b0;
    assign data[3807] = 16'b0;
    assign data[3808] = 16'b0;
    assign data[3809] = 16'b0;
    assign data[3810] = 16'b0;
    assign data[3811] = 16'b0;
    assign data[3812] = ~16'b0;
    assign data[3813] = ~16'b0;
    assign data[3814] = ~16'b0;
    assign data[3815] = ~16'b0;
    assign data[3816] = ~16'b0;
    assign data[3817] = ~16'b0;
    assign data[3818] = ~16'b0;
    assign data[3819] = ~16'b0;
    assign data[3820] = 16'b0;
    assign data[3821] = 16'b0;
    assign data[3822] = ~16'b0;
    assign data[3823] = ~16'b0;
    assign data[3824] = ~16'b0;
    assign data[3825] = ~16'b0;
    assign data[3826] = ~16'b0;
    assign data[3827] = ~16'b0;
    assign data[3828] = ~16'b0;
    assign data[3829] = ~16'b0;
    assign data[3830] = 16'b0;
    assign data[3831] = 16'b0;
    assign data[3832] = ~16'b0;
    assign data[3833] = ~16'b0;
    assign data[3834] = ~16'b0;
    assign data[3835] = ~16'b0;
    assign data[3836] = ~16'b0;
    assign data[3837] = ~16'b0;
    assign data[3838] = ~16'b0;
    assign data[3839] = ~16'b0;
    assign data[3840] = 16'b0;
    assign data[3841] = 16'b0;
    assign data[3842] = ~16'b0;
    assign data[3843] = ~16'b0;
    assign data[3844] = ~16'b0;
    assign data[3845] = ~16'b0;
    assign data[3846] = ~16'b0;
    assign data[3847] = ~16'b0;
    assign data[3848] = ~16'b0;
    assign data[3849] = ~16'b0;
    assign data[3850] = 16'b0;
    assign data[3851] = 16'b0;
    assign data[3852] = ~16'b0;
    assign data[3853] = ~16'b0;
    assign data[3854] = ~16'b0;
    assign data[3855] = ~16'b0;
    assign data[3856] = ~16'b0;
    assign data[3857] = ~16'b0;
    assign data[3858] = ~16'b0;
    assign data[3859] = ~16'b0;
    assign data[3860] = 16'b0;
    assign data[3861] = 16'b0;
    assign data[3862] = ~16'b0;
    assign data[3863] = ~16'b0;
    assign data[3864] = ~16'b0;
    assign data[3865] = ~16'b0;
    assign data[3866] = ~16'b0;
    assign data[3867] = ~16'b0;
    assign data[3868] = ~16'b0;
    assign data[3869] = ~16'b0;
    assign data[3870] = 16'b0;
    assign data[3871] = 16'b0;
    assign data[3872] = ~16'b0;
    assign data[3873] = ~16'b0;
    assign data[3874] = ~16'b0;
    assign data[3875] = ~16'b0;
    assign data[3876] = ~16'b0;
    assign data[3877] = ~16'b0;
    assign data[3878] = ~16'b0;
    assign data[3879] = ~16'b0;
    assign data[3880] = 16'b0;
    assign data[3881] = 16'b0;
    assign data[3882] = ~16'b0;
    assign data[3883] = ~16'b0;
    assign data[3884] = ~16'b0;
    assign data[3885] = ~16'b0;
    assign data[3886] = ~16'b0;
    assign data[3887] = ~16'b0;
    assign data[3888] = ~16'b0;
    assign data[3889] = ~16'b0;
    assign data[3890] = 16'b0;
    assign data[3891] = 16'b0;
    assign data[3892] = ~16'b0;
    assign data[3893] = ~16'b0;
    assign data[3894] = ~16'b0;
    assign data[3895] = ~16'b0;
    assign data[3896] = ~16'b0;
    assign data[3897] = ~16'b0;
    assign data[3898] = ~16'b0;
    assign data[3899] = ~16'b0;
    assign data[3900] = 16'b0;
    assign data[3901] = 16'b0;
    assign data[3902] = ~16'b0;
    assign data[3903] = ~16'b0;
    assign data[3904] = ~16'b0;
    assign data[3905] = ~16'b0;
    assign data[3906] = ~16'b0;
    assign data[3907] = ~16'b0;
    assign data[3908] = ~16'b0;
    assign data[3909] = ~16'b0;
    assign data[3910] = 16'b0;
    assign data[3911] = 16'b0;
    assign data[3912] = ~16'b0;
    assign data[3913] = ~16'b0;
    assign data[3914] = ~16'b0;
    assign data[3915] = ~16'b0;
    assign data[3916] = ~16'b0;
    assign data[3917] = ~16'b0;
    assign data[3918] = ~16'b0;
    assign data[3919] = ~16'b0;
    assign data[3920] = 16'b0;
    assign data[3921] = 16'b0;
    assign data[3922] = ~16'b0;
    assign data[3923] = ~16'b0;
    assign data[3924] = ~16'b0;
    assign data[3925] = ~16'b0;
    assign data[3926] = ~16'b0;
    assign data[3927] = ~16'b0;
    assign data[3928] = ~16'b0;
    assign data[3929] = ~16'b0;
    assign data[3930] = 16'b0;
    assign data[3931] = 16'b0;
    assign data[3932] = ~16'b0;
    assign data[3933] = ~16'b0;
    assign data[3934] = ~16'b0;
    assign data[3935] = ~16'b0;
    assign data[3936] = ~16'b0;
    assign data[3937] = ~16'b0;
    assign data[3938] = ~16'b0;
    assign data[3939] = ~16'b0;
    assign data[3940] = 16'b0;
    assign data[3941] = 16'b0;
    assign data[3942] = ~16'b0;
    assign data[3943] = ~16'b0;
    assign data[3944] = ~16'b0;
    assign data[3945] = ~16'b0;
    assign data[3946] = ~16'b0;
    assign data[3947] = ~16'b0;
    assign data[3948] = ~16'b0;
    assign data[3949] = ~16'b0;
    assign data[3950] = 16'b0;
    assign data[3951] = 16'b0;
    assign data[3952] = ~16'b0;
    assign data[3953] = ~16'b0;
    assign data[3954] = ~16'b0;
    assign data[3955] = ~16'b0;
    assign data[3956] = ~16'b0;
    assign data[3957] = ~16'b0;
    assign data[3958] = ~16'b0;
    assign data[3959] = ~16'b0;
    assign data[3960] = 16'b0;
    assign data[3961] = 16'b0;
    assign data[3962] = ~16'b0;
    assign data[3963] = ~16'b0;
    assign data[3964] = ~16'b0;
    assign data[3965] = ~16'b0;
    assign data[3966] = ~16'b0;
    assign data[3967] = ~16'b0;
    assign data[3968] = ~16'b0;
    assign data[3969] = ~16'b0;
    assign data[3970] = 16'b0;
    assign data[3971] = 16'b0;
    assign data[3972] = ~16'b0;
    assign data[3973] = ~16'b0;
    assign data[3974] = ~16'b0;
    assign data[3975] = ~16'b0;
    assign data[3976] = ~16'b0;
    assign data[3977] = ~16'b0;
    assign data[3978] = ~16'b0;
    assign data[3979] = ~16'b0;
    assign data[3980] = 16'b0;
    assign data[3981] = 16'b0;
    assign data[3982] = ~16'b0;
    assign data[3983] = ~16'b0;
    assign data[3984] = ~16'b0;
    assign data[3985] = ~16'b0;
    assign data[3986] = ~16'b0;
    assign data[3987] = ~16'b0;
    assign data[3988] = ~16'b0;
    assign data[3989] = ~16'b0;
    assign data[3990] = 16'b0;
    assign data[3991] = 16'b0;
    assign data[3992] = ~16'b0;
    assign data[3993] = ~16'b0;
    assign data[3994] = ~16'b0;
    assign data[3995] = ~16'b0;
    assign data[3996] = ~16'b0;
    assign data[3997] = ~16'b0;
    assign data[3998] = ~16'b0;
    assign data[3999] = ~16'b0;
    assign data[4000] = 16'b0;
    assign data[4001] = 16'b0;
    assign data[4002] = ~16'b0;
    assign data[4003] = ~16'b0;
    assign data[4004] = ~16'b0;
    assign data[4005] = ~16'b0;
    assign data[4006] = ~16'b0;
    assign data[4007] = ~16'b0;
    assign data[4008] = ~16'b0;
    assign data[4009] = ~16'b0;
    assign data[4010] = 16'b0;
    assign data[4011] = 16'b0;
    assign data[4012] = ~16'b0;
    assign data[4013] = ~16'b0;
    assign data[4014] = ~16'b0;
    assign data[4015] = ~16'b0;
    assign data[4016] = ~16'b0;
    assign data[4017] = ~16'b0;
    assign data[4018] = ~16'b0;
    assign data[4019] = ~16'b0;
    assign data[4020] = 16'b0;
    assign data[4021] = 16'b0;
    assign data[4022] = ~16'b0;
    assign data[4023] = ~16'b0;
    assign data[4024] = ~16'b0;
    assign data[4025] = ~16'b0;
    assign data[4026] = ~16'b0;
    assign data[4027] = ~16'b0;
    assign data[4028] = ~16'b0;
    assign data[4029] = ~16'b0;
    assign data[4030] = 16'b0;
    assign data[4031] = 16'b0;
    assign data[4032] = ~16'b0;
    assign data[4033] = ~16'b0;
    assign data[4034] = ~16'b0;
    assign data[4035] = ~16'b0;
    assign data[4036] = ~16'b0;
    assign data[4037] = ~16'b0;
    assign data[4038] = ~16'b0;
    assign data[4039] = ~16'b0;
    assign data[4040] = 16'b0;
    assign data[4041] = 16'b0;
    assign data[4042] = ~16'b0;
    assign data[4043] = ~16'b0;
    assign data[4044] = ~16'b0;
    assign data[4045] = ~16'b0;
    assign data[4046] = ~16'b0;
    assign data[4047] = ~16'b0;
    assign data[4048] = ~16'b0;
    assign data[4049] = ~16'b0;
    assign data[4050] = 16'b0;
    assign data[4051] = 16'b0;
    assign data[4052] = ~16'b0;
    assign data[4053] = ~16'b0;
    assign data[4054] = ~16'b0;
    assign data[4055] = ~16'b0;
    assign data[4056] = ~16'b0;
    assign data[4057] = ~16'b0;
    assign data[4058] = ~16'b0;
    assign data[4059] = ~16'b0;
    assign data[4060] = 16'b0;
    assign data[4061] = 16'b0;
    assign data[4062] = ~16'b0;
    assign data[4063] = ~16'b0;
    assign data[4064] = ~16'b0;
    assign data[4065] = ~16'b0;
    assign data[4066] = ~16'b0;
    assign data[4067] = ~16'b0;
    assign data[4068] = ~16'b0;
    assign data[4069] = ~16'b0;
    assign data[4070] = 16'b0;
    assign data[4071] = 16'b0;
    assign data[4072] = ~16'b0;
    assign data[4073] = ~16'b0;
    assign data[4074] = ~16'b0;
    assign data[4075] = ~16'b0;
    assign data[4076] = ~16'b0;
    assign data[4077] = ~16'b0;
    assign data[4078] = ~16'b0;
    assign data[4079] = ~16'b0;
    assign data[4080] = 16'b0;
    assign data[4081] = 16'b0;
    assign data[4082] = ~16'b0;
    assign data[4083] = ~16'b0;
    assign data[4084] = ~16'b0;
    assign data[4085] = ~16'b0;
    assign data[4086] = ~16'b0;
    assign data[4087] = ~16'b0;
    assign data[4088] = ~16'b0;
    assign data[4089] = ~16'b0;
    assign data[4090] = 16'b0;
    assign data[4091] = 16'b0;
    assign data[4092] = ~16'b0;
    assign data[4093] = ~16'b0;
    assign data[4094] = ~16'b0;
    assign data[4095] = ~16'b0;
    assign data[4096] = ~16'b0;
    assign data[4097] = ~16'b0;
    assign data[4098] = ~16'b0;
    assign data[4099] = ~16'b0;
    assign data[4100] = 16'b0;
    assign data[4101] = 16'b0;
    assign data[4102] = ~16'b0;
    assign data[4103] = ~16'b0;
    assign data[4104] = ~16'b0;
    assign data[4105] = ~16'b0;
    assign data[4106] = ~16'b0;
    assign data[4107] = ~16'b0;
    assign data[4108] = ~16'b0;
    assign data[4109] = ~16'b0;
    assign data[4110] = 16'b0;
    assign data[4111] = 16'b0;
    assign data[4112] = ~16'b0;
    assign data[4113] = ~16'b0;
    assign data[4114] = ~16'b0;
    assign data[4115] = ~16'b0;
    assign data[4116] = ~16'b0;
    assign data[4117] = ~16'b0;
    assign data[4118] = ~16'b0;
    assign data[4119] = ~16'b0;
    assign data[4120] = 16'b0;
    assign data[4121] = 16'b0;
    assign data[4122] = ~16'b0;
    assign data[4123] = ~16'b0;
    assign data[4124] = ~16'b0;
    assign data[4125] = ~16'b0;
    assign data[4126] = ~16'b0;
    assign data[4127] = ~16'b0;
    assign data[4128] = ~16'b0;
    assign data[4129] = ~16'b0;
    assign data[4130] = 16'b0;
    assign data[4131] = 16'b0;
    assign data[4132] = ~16'b0;
    assign data[4133] = ~16'b0;
    assign data[4134] = ~16'b0;
    assign data[4135] = ~16'b0;
    assign data[4136] = ~16'b0;
    assign data[4137] = ~16'b0;
    assign data[4138] = ~16'b0;
    assign data[4139] = ~16'b0;
    assign data[4140] = 16'b0;
    assign data[4141] = 16'b0;
    assign data[4142] = ~16'b0;
    assign data[4143] = ~16'b0;
    assign data[4144] = ~16'b0;
    assign data[4145] = ~16'b0;
    assign data[4146] = ~16'b0;
    assign data[4147] = ~16'b0;
    assign data[4148] = ~16'b0;
    assign data[4149] = ~16'b0;
    assign data[4150] = 16'b0;
    assign data[4151] = 16'b0;
    assign data[4152] = 16'b0;
    assign data[4153] = 16'b0;
    assign data[4154] = 16'b0;
    assign data[4155] = 16'b0;
    assign data[4156] = 16'b0;
    assign data[4157] = 16'b0;
    assign data[4158] = 16'b0;
    assign data[4159] = 16'b0;
    assign data[4160] = 16'b0;
    assign data[4161] = 16'b0;
    assign data[4162] = 16'b0;
    assign data[4163] = 16'b0;
    assign data[4164] = 16'b0;
    assign data[4165] = 16'b0;
    assign data[4166] = 16'b0;
    assign data[4167] = 16'b0;
    assign data[4168] = 16'b0;
    assign data[4169] = 16'b0;
    assign data[4170] = ~16'b0;
    assign data[4171] = ~16'b0;
    assign data[4172] = ~16'b0;
    assign data[4173] = ~16'b0;
    assign data[4174] = ~16'b0;
    assign data[4175] = ~16'b0;
    assign data[4176] = ~16'b0;
    assign data[4177] = ~16'b0;
    assign data[4178] = ~16'b0;
    assign data[4179] = ~16'b0;
    assign data[4180] = ~16'b0;
    assign data[4181] = ~16'b0;
    assign data[4182] = ~16'b0;
    assign data[4183] = ~16'b0;
    assign data[4184] = ~16'b0;
    assign data[4185] = ~16'b0;
    assign data[4186] = ~16'b0;
    assign data[4187] = ~16'b0;
    assign data[4188] = ~16'b0;
    assign data[4189] = ~16'b0;
    assign data[4190] = ~16'b0;
    assign data[4191] = ~16'b0;
    assign data[4192] = ~16'b0;
    assign data[4193] = ~16'b0;
    assign data[4194] = ~16'b0;
    assign data[4195] = ~16'b0;
    assign data[4196] = ~16'b0;
    assign data[4197] = ~16'b0;
    assign data[4198] = ~16'b0;
    assign data[4199] = ~16'b0;
    assign data[4200] = ~16'b0;
    assign data[4201] = ~16'b0;
    assign data[4202] = ~16'b0;
    assign data[4203] = ~16'b0;
    assign data[4204] = ~16'b0;
    assign data[4205] = ~16'b0;
    assign data[4206] = ~16'b0;
    assign data[4207] = ~16'b0;
    assign data[4208] = ~16'b0;
    assign data[4209] = ~16'b0;
    assign data[4210] = ~16'b0;
    assign data[4211] = ~16'b0;
    assign data[4212] = ~16'b0;
    assign data[4213] = ~16'b0;
    assign data[4214] = ~16'b0;
    assign data[4215] = ~16'b0;
    assign data[4216] = ~16'b0;
    assign data[4217] = ~16'b0;
    assign data[4218] = ~16'b0;
    assign data[4219] = ~16'b0;
    assign data[4220] = ~16'b0;
    assign data[4221] = ~16'b0;
    assign data[4222] = ~16'b0;
    assign data[4223] = ~16'b0;
    assign data[4224] = ~16'b0;
    assign data[4225] = ~16'b0;
    assign data[4226] = ~16'b0;
    assign data[4227] = ~16'b0;
    assign data[4228] = ~16'b0;
    assign data[4229] = ~16'b0;
    assign data[4230] = ~16'b0;
    assign data[4231] = ~16'b0;
    assign data[4232] = ~16'b0;
    assign data[4233] = ~16'b0;
    assign data[4234] = ~16'b0;
    assign data[4235] = ~16'b0;
    assign data[4236] = ~16'b0;
    assign data[4237] = ~16'b0;
    assign data[4238] = ~16'b0;
    assign data[4239] = ~16'b0;
    assign data[4240] = ~16'b0;
    assign data[4241] = ~16'b0;
    assign data[4242] = ~16'b0;
    assign data[4243] = ~16'b0;
    assign data[4244] = ~16'b0;
    assign data[4245] = ~16'b0;
    assign data[4246] = ~16'b0;
    assign data[4247] = ~16'b0;
    assign data[4248] = ~16'b0;
    assign data[4249] = ~16'b0;
    assign data[4250] = ~16'b0;
    assign data[4251] = ~16'b0;
    assign data[4252] = ~16'b0;
    assign data[4253] = ~16'b0;
    assign data[4254] = ~16'b0;
    assign data[4255] = ~16'b0;
    assign data[4256] = ~16'b0;
    assign data[4257] = ~16'b0;
    assign data[4258] = ~16'b0;
    assign data[4259] = ~16'b0;
    assign data[4260] = ~16'b0;
    assign data[4261] = ~16'b0;
    assign data[4262] = ~16'b0;
    assign data[4263] = ~16'b0;
    assign data[4264] = ~16'b0;
    assign data[4265] = ~16'b0;
    assign data[4266] = ~16'b0;
    assign data[4267] = ~16'b0;
    assign data[4268] = ~16'b0;
    assign data[4269] = ~16'b0;
    assign data[4270] = 16'b0;
    assign data[4271] = 16'b0;
    assign data[4272] = 16'b0;
    assign data[4273] = 16'b0;
    assign data[4274] = 16'b0;
    assign data[4275] = 16'b0;
    assign data[4276] = 16'b0;
    assign data[4277] = 16'b0;
    assign data[4278] = 16'b0;
    assign data[4279] = 16'b0;
    assign data[4280] = 16'b0;
    assign data[4281] = 16'b0;
    assign data[4282] = 16'b0;
    assign data[4283] = 16'b0;
    assign data[4284] = 16'b0;
    assign data[4285] = 16'b0;
    assign data[4286] = 16'b0;
    assign data[4287] = 16'b0;
    assign data[4288] = 16'b0;
    assign data[4289] = 16'b0;
    assign data[4290] = 16'b0;
    assign data[4291] = 16'b0;
    assign data[4292] = ~16'b0;
    assign data[4293] = ~16'b0;
    assign data[4294] = ~16'b0;
    assign data[4295] = ~16'b0;
    assign data[4296] = ~16'b0;
    assign data[4297] = ~16'b0;
    assign data[4298] = ~16'b0;
    assign data[4299] = ~16'b0;
    assign data[4300] = 16'b0;
    assign data[4301] = 16'b0;
    assign data[4302] = ~16'b0;
    assign data[4303] = ~16'b0;
    assign data[4304] = ~16'b0;
    assign data[4305] = ~16'b0;
    assign data[4306] = ~16'b0;
    assign data[4307] = ~16'b0;
    assign data[4308] = ~16'b0;
    assign data[4309] = ~16'b0;
    assign data[4310] = 16'b0;
    assign data[4311] = 16'b0;
    assign data[4312] = ~16'b0;
    assign data[4313] = ~16'b0;
    assign data[4314] = ~16'b0;
    assign data[4315] = ~16'b0;
    assign data[4316] = ~16'b0;
    assign data[4317] = ~16'b0;
    assign data[4318] = ~16'b0;
    assign data[4319] = ~16'b0;
    assign data[4320] = 16'b0;
    assign data[4321] = 16'b0;
    assign data[4322] = ~16'b0;
    assign data[4323] = ~16'b0;
    assign data[4324] = ~16'b0;
    assign data[4325] = ~16'b0;
    assign data[4326] = ~16'b0;
    assign data[4327] = ~16'b0;
    assign data[4328] = ~16'b0;
    assign data[4329] = ~16'b0;
    assign data[4330] = 16'b0;
    assign data[4331] = 16'b0;
    assign data[4332] = ~16'b0;
    assign data[4333] = ~16'b0;
    assign data[4334] = ~16'b0;
    assign data[4335] = ~16'b0;
    assign data[4336] = ~16'b0;
    assign data[4337] = ~16'b0;
    assign data[4338] = ~16'b0;
    assign data[4339] = ~16'b0;
    assign data[4340] = 16'b0;
    assign data[4341] = 16'b0;
    assign data[4342] = ~16'b0;
    assign data[4343] = ~16'b0;
    assign data[4344] = ~16'b0;
    assign data[4345] = ~16'b0;
    assign data[4346] = ~16'b0;
    assign data[4347] = ~16'b0;
    assign data[4348] = ~16'b0;
    assign data[4349] = ~16'b0;
    assign data[4350] = 16'b0;
    assign data[4351] = 16'b0;
    assign data[4352] = ~16'b0;
    assign data[4353] = ~16'b0;
    assign data[4354] = ~16'b0;
    assign data[4355] = ~16'b0;
    assign data[4356] = ~16'b0;
    assign data[4357] = ~16'b0;
    assign data[4358] = ~16'b0;
    assign data[4359] = ~16'b0;
    assign data[4360] = 16'b0;
    assign data[4361] = 16'b0;
    assign data[4362] = ~16'b0;
    assign data[4363] = ~16'b0;
    assign data[4364] = ~16'b0;
    assign data[4365] = ~16'b0;
    assign data[4366] = ~16'b0;
    assign data[4367] = ~16'b0;
    assign data[4368] = ~16'b0;
    assign data[4369] = ~16'b0;
    assign data[4370] = 16'b0;
    assign data[4371] = 16'b0;
    assign data[4372] = ~16'b0;
    assign data[4373] = ~16'b0;
    assign data[4374] = ~16'b0;
    assign data[4375] = ~16'b0;
    assign data[4376] = ~16'b0;
    assign data[4377] = ~16'b0;
    assign data[4378] = ~16'b0;
    assign data[4379] = ~16'b0;
    assign data[4380] = 16'b0;
    assign data[4381] = 16'b0;
    assign data[4382] = ~16'b0;
    assign data[4383] = ~16'b0;
    assign data[4384] = ~16'b0;
    assign data[4385] = ~16'b0;
    assign data[4386] = ~16'b0;
    assign data[4387] = ~16'b0;
    assign data[4388] = ~16'b0;
    assign data[4389] = ~16'b0;
    assign data[4390] = 16'b0;
    assign data[4391] = 16'b0;
    assign data[4392] = ~16'b0;
    assign data[4393] = ~16'b0;
    assign data[4394] = ~16'b0;
    assign data[4395] = ~16'b0;
    assign data[4396] = ~16'b0;
    assign data[4397] = ~16'b0;
    assign data[4398] = ~16'b0;
    assign data[4399] = ~16'b0;
    assign data[4400] = 16'b0;
    assign data[4401] = 16'b0;
    assign data[4402] = ~16'b0;
    assign data[4403] = ~16'b0;
    assign data[4404] = ~16'b0;
    assign data[4405] = ~16'b0;
    assign data[4406] = ~16'b0;
    assign data[4407] = ~16'b0;
    assign data[4408] = ~16'b0;
    assign data[4409] = ~16'b0;
    assign data[4410] = 16'b0;
    assign data[4411] = 16'b0;
    assign data[4412] = ~16'b0;
    assign data[4413] = ~16'b0;
    assign data[4414] = ~16'b0;
    assign data[4415] = ~16'b0;
    assign data[4416] = ~16'b0;
    assign data[4417] = ~16'b0;
    assign data[4418] = ~16'b0;
    assign data[4419] = ~16'b0;
    assign data[4420] = 16'b0;
    assign data[4421] = 16'b0;
    assign data[4422] = ~16'b0;
    assign data[4423] = ~16'b0;
    assign data[4424] = ~16'b0;
    assign data[4425] = ~16'b0;
    assign data[4426] = ~16'b0;
    assign data[4427] = ~16'b0;
    assign data[4428] = ~16'b0;
    assign data[4429] = ~16'b0;
    assign data[4430] = 16'b0;
    assign data[4431] = 16'b0;
    assign data[4432] = ~16'b0;
    assign data[4433] = ~16'b0;
    assign data[4434] = ~16'b0;
    assign data[4435] = ~16'b0;
    assign data[4436] = ~16'b0;
    assign data[4437] = ~16'b0;
    assign data[4438] = ~16'b0;
    assign data[4439] = ~16'b0;
    assign data[4440] = 16'b0;
    assign data[4441] = 16'b0;
    assign data[4442] = ~16'b0;
    assign data[4443] = ~16'b0;
    assign data[4444] = ~16'b0;
    assign data[4445] = ~16'b0;
    assign data[4446] = ~16'b0;
    assign data[4447] = ~16'b0;
    assign data[4448] = ~16'b0;
    assign data[4449] = ~16'b0;
    assign data[4450] = 16'b0;
    assign data[4451] = 16'b0;
    assign data[4452] = ~16'b0;
    assign data[4453] = ~16'b0;
    assign data[4454] = ~16'b0;
    assign data[4455] = ~16'b0;
    assign data[4456] = ~16'b0;
    assign data[4457] = ~16'b0;
    assign data[4458] = ~16'b0;
    assign data[4459] = ~16'b0;
    assign data[4460] = 16'b0;
    assign data[4461] = 16'b0;
    assign data[4462] = ~16'b0;
    assign data[4463] = ~16'b0;
    assign data[4464] = ~16'b0;
    assign data[4465] = ~16'b0;
    assign data[4466] = ~16'b0;
    assign data[4467] = ~16'b0;
    assign data[4468] = ~16'b0;
    assign data[4469] = ~16'b0;
    assign data[4470] = 16'b0;
    assign data[4471] = 16'b0;
    assign data[4472] = ~16'b0;
    assign data[4473] = ~16'b0;
    assign data[4474] = ~16'b0;
    assign data[4475] = ~16'b0;
    assign data[4476] = ~16'b0;
    assign data[4477] = ~16'b0;
    assign data[4478] = ~16'b0;
    assign data[4479] = ~16'b0;
    assign data[4480] = 16'b0;
    assign data[4481] = 16'b0;
    assign data[4482] = ~16'b0;
    assign data[4483] = ~16'b0;
    assign data[4484] = ~16'b0;
    assign data[4485] = ~16'b0;
    assign data[4486] = ~16'b0;
    assign data[4487] = ~16'b0;
    assign data[4488] = ~16'b0;
    assign data[4489] = ~16'b0;
    assign data[4490] = 16'b0;
    assign data[4491] = 16'b0;
    assign data[4492] = ~16'b0;
    assign data[4493] = ~16'b0;
    assign data[4494] = ~16'b0;
    assign data[4495] = ~16'b0;
    assign data[4496] = ~16'b0;
    assign data[4497] = ~16'b0;
    assign data[4498] = ~16'b0;
    assign data[4499] = ~16'b0;
    assign data[4500] = 16'b0;
    assign data[4501] = 16'b0;
    assign data[4502] = ~16'b0;
    assign data[4503] = ~16'b0;
    assign data[4504] = ~16'b0;
    assign data[4505] = ~16'b0;
    assign data[4506] = ~16'b0;
    assign data[4507] = ~16'b0;
    assign data[4508] = ~16'b0;
    assign data[4509] = ~16'b0;
    assign data[4510] = 16'b0;
    assign data[4511] = 16'b0;
    assign data[4512] = ~16'b0;
    assign data[4513] = ~16'b0;
    assign data[4514] = ~16'b0;
    assign data[4515] = ~16'b0;
    assign data[4516] = ~16'b0;
    assign data[4517] = ~16'b0;
    assign data[4518] = ~16'b0;
    assign data[4519] = ~16'b0;
    assign data[4520] = 16'b0;
    assign data[4521] = 16'b0;
    assign data[4522] = ~16'b0;
    assign data[4523] = ~16'b0;
    assign data[4524] = ~16'b0;
    assign data[4525] = ~16'b0;
    assign data[4526] = ~16'b0;
    assign data[4527] = ~16'b0;
    assign data[4528] = ~16'b0;
    assign data[4529] = ~16'b0;
    assign data[4530] = 16'b0;
    assign data[4531] = 16'b0;
    assign data[4532] = ~16'b0;
    assign data[4533] = ~16'b0;
    assign data[4534] = ~16'b0;
    assign data[4535] = ~16'b0;
    assign data[4536] = ~16'b0;
    assign data[4537] = ~16'b0;
    assign data[4538] = ~16'b0;
    assign data[4539] = ~16'b0;
    assign data[4540] = 16'b0;
    assign data[4541] = 16'b0;
    assign data[4542] = ~16'b0;
    assign data[4543] = ~16'b0;
    assign data[4544] = ~16'b0;
    assign data[4545] = ~16'b0;
    assign data[4546] = ~16'b0;
    assign data[4547] = ~16'b0;
    assign data[4548] = ~16'b0;
    assign data[4549] = ~16'b0;
    assign data[4550] = 16'b0;
    assign data[4551] = 16'b0;
    assign data[4552] = ~16'b0;
    assign data[4553] = ~16'b0;
    assign data[4554] = ~16'b0;
    assign data[4555] = ~16'b0;
    assign data[4556] = ~16'b0;
    assign data[4557] = ~16'b0;
    assign data[4558] = ~16'b0;
    assign data[4559] = ~16'b0;
    assign data[4560] = 16'b0;
    assign data[4561] = 16'b0;
    assign data[4562] = ~16'b0;
    assign data[4563] = ~16'b0;
    assign data[4564] = ~16'b0;
    assign data[4565] = ~16'b0;
    assign data[4566] = ~16'b0;
    assign data[4567] = ~16'b0;
    assign data[4568] = ~16'b0;
    assign data[4569] = ~16'b0;
    assign data[4570] = 16'b0;
    assign data[4571] = 16'b0;
    assign data[4572] = ~16'b0;
    assign data[4573] = ~16'b0;
    assign data[4574] = ~16'b0;
    assign data[4575] = ~16'b0;
    assign data[4576] = ~16'b0;
    assign data[4577] = ~16'b0;
    assign data[4578] = ~16'b0;
    assign data[4579] = ~16'b0;
    assign data[4580] = 16'b0;
    assign data[4581] = 16'b0;
    assign data[4582] = ~16'b0;
    assign data[4583] = ~16'b0;
    assign data[4584] = ~16'b0;
    assign data[4585] = ~16'b0;
    assign data[4586] = ~16'b0;
    assign data[4587] = ~16'b0;
    assign data[4588] = ~16'b0;
    assign data[4589] = ~16'b0;
    assign data[4590] = 16'b0;
    assign data[4591] = 16'b0;
    assign data[4592] = ~16'b0;
    assign data[4593] = ~16'b0;
    assign data[4594] = ~16'b0;
    assign data[4595] = ~16'b0;
    assign data[4596] = ~16'b0;
    assign data[4597] = ~16'b0;
    assign data[4598] = ~16'b0;
    assign data[4599] = ~16'b0;
    assign data[4600] = 16'b0;
    assign data[4601] = 16'b0;
    assign data[4602] = ~16'b0;
    assign data[4603] = ~16'b0;
    assign data[4604] = ~16'b0;
    assign data[4605] = ~16'b0;
    assign data[4606] = ~16'b0;
    assign data[4607] = ~16'b0;
    assign data[4608] = ~16'b0;
    assign data[4609] = ~16'b0;
    assign data[4610] = 16'b0;
    assign data[4611] = 16'b0;
    assign data[4612] = ~16'b0;
    assign data[4613] = ~16'b0;
    assign data[4614] = ~16'b0;
    assign data[4615] = ~16'b0;
    assign data[4616] = ~16'b0;
    assign data[4617] = ~16'b0;
    assign data[4618] = ~16'b0;
    assign data[4619] = ~16'b0;
    assign data[4620] = 16'b0;
    assign data[4621] = 16'b0;
    assign data[4622] = ~16'b0;
    assign data[4623] = ~16'b0;
    assign data[4624] = ~16'b0;
    assign data[4625] = ~16'b0;
    assign data[4626] = ~16'b0;
    assign data[4627] = ~16'b0;
    assign data[4628] = ~16'b0;
    assign data[4629] = ~16'b0;
    assign data[4630] = 16'b0;
    assign data[4631] = 16'b0;
    assign data[4632] = ~16'b0;
    assign data[4633] = ~16'b0;
    assign data[4634] = ~16'b0;
    assign data[4635] = ~16'b0;
    assign data[4636] = ~16'b0;
    assign data[4637] = ~16'b0;
    assign data[4638] = ~16'b0;
    assign data[4639] = ~16'b0;
    assign data[4640] = 16'b0;
    assign data[4641] = 16'b0;
    assign data[4642] = ~16'b0;
    assign data[4643] = ~16'b0;
    assign data[4644] = ~16'b0;
    assign data[4645] = ~16'b0;
    assign data[4646] = ~16'b0;
    assign data[4647] = ~16'b0;
    assign data[4648] = ~16'b0;
    assign data[4649] = ~16'b0;
    assign data[4650] = 16'b0;
    assign data[4651] = 16'b0;
    assign data[4652] = 16'b0;
    assign data[4653] = 16'b0;
    assign data[4654] = 16'b0;
    assign data[4655] = 16'b0;
    assign data[4656] = 16'b0;
    assign data[4657] = 16'b0;
    assign data[4658] = 16'b0;
    assign data[4659] = 16'b0;
    assign data[4660] = 16'b0;
    assign data[4661] = 16'b0;
    assign data[4662] = 16'b0;
    assign data[4663] = 16'b0;
    assign data[4664] = 16'b0;
    assign data[4665] = 16'b0;
    assign data[4666] = 16'b0;
    assign data[4667] = 16'b0;
    assign data[4668] = 16'b0;
    assign data[4669] = 16'b0;
    assign data[4670] = ~16'b0;
    assign data[4671] = ~16'b0;
    assign data[4672] = ~16'b0;
    assign data[4673] = ~16'b0;
    assign data[4674] = ~16'b0;
    assign data[4675] = ~16'b0;
    assign data[4676] = ~16'b0;
    assign data[4677] = ~16'b0;
    assign data[4678] = ~16'b0;
    assign data[4679] = ~16'b0;
    assign data[4680] = ~16'b0;
    assign data[4681] = ~16'b0;
    assign data[4682] = ~16'b0;
    assign data[4683] = ~16'b0;
    assign data[4684] = ~16'b0;
    assign data[4685] = ~16'b0;
    assign data[4686] = ~16'b0;
    assign data[4687] = ~16'b0;
    assign data[4688] = ~16'b0;
    assign data[4689] = ~16'b0;
    assign data[4690] = ~16'b0;
    assign data[4691] = ~16'b0;
    assign data[4692] = ~16'b0;
    assign data[4693] = ~16'b0;
    assign data[4694] = ~16'b0;
    assign data[4695] = ~16'b0;
    assign data[4696] = ~16'b0;
    assign data[4697] = ~16'b0;
    assign data[4698] = ~16'b0;
    assign data[4699] = ~16'b0;
    assign data[4700] = ~16'b0;
    assign data[4701] = ~16'b0;
    assign data[4702] = ~16'b0;
    assign data[4703] = ~16'b0;
    assign data[4704] = ~16'b0;
    assign data[4705] = ~16'b0;
    assign data[4706] = ~16'b0;
    assign data[4707] = ~16'b0;
    assign data[4708] = ~16'b0;
    assign data[4709] = ~16'b0;
    assign data[4710] = ~16'b0;
    assign data[4711] = ~16'b0;
    assign data[4712] = ~16'b0;
    assign data[4713] = ~16'b0;
    assign data[4714] = ~16'b0;
    assign data[4715] = ~16'b0;
    assign data[4716] = ~16'b0;
    assign data[4717] = ~16'b0;
    assign data[4718] = ~16'b0;
    assign data[4719] = ~16'b0;
    assign data[4720] = ~16'b0;
    assign data[4721] = ~16'b0;
    assign data[4722] = ~16'b0;
    assign data[4723] = ~16'b0;
    assign data[4724] = ~16'b0;
    assign data[4725] = ~16'b0;
    assign data[4726] = ~16'b0;
    assign data[4727] = ~16'b0;
    assign data[4728] = ~16'b0;
    assign data[4729] = ~16'b0;
    assign data[4730] = ~16'b0;
    assign data[4731] = ~16'b0;
    assign data[4732] = ~16'b0;
    assign data[4733] = ~16'b0;
    assign data[4734] = ~16'b0;
    assign data[4735] = ~16'b0;
    assign data[4736] = ~16'b0;
    assign data[4737] = ~16'b0;
    assign data[4738] = ~16'b0;
    assign data[4739] = ~16'b0;
    assign data[4740] = ~16'b0;
    assign data[4741] = ~16'b0;
    assign data[4742] = ~16'b0;
    assign data[4743] = ~16'b0;
    assign data[4744] = ~16'b0;
    assign data[4745] = ~16'b0;
    assign data[4746] = ~16'b0;
    assign data[4747] = ~16'b0;
    assign data[4748] = ~16'b0;
    assign data[4749] = ~16'b0;
    assign data[4750] = ~16'b0;
    assign data[4751] = ~16'b0;
    assign data[4752] = ~16'b0;
    assign data[4753] = ~16'b0;
    assign data[4754] = ~16'b0;
    assign data[4755] = ~16'b0;
    assign data[4756] = ~16'b0;
    assign data[4757] = ~16'b0;
    assign data[4758] = ~16'b0;
    assign data[4759] = ~16'b0;
    assign data[4760] = ~16'b0;
    assign data[4761] = ~16'b0;
    assign data[4762] = ~16'b0;
    assign data[4763] = ~16'b0;
    assign data[4764] = ~16'b0;
    assign data[4765] = ~16'b0;
    assign data[4766] = ~16'b0;
    assign data[4767] = ~16'b0;
    assign data[4768] = ~16'b0;
    assign data[4769] = ~16'b0;
    assign data[4770] = ~16'b0;
    assign data[4771] = ~16'b0;
    assign data[4772] = ~16'b0;
    assign data[4773] = ~16'b0;
    assign data[4774] = ~16'b0;
    assign data[4775] = ~16'b0;
    assign data[4776] = ~16'b0;
    assign data[4777] = ~16'b0;
    assign data[4778] = ~16'b0;
    assign data[4779] = ~16'b0;
    assign data[4780] = ~16'b0;
    assign data[4781] = ~16'b0;
    assign data[4782] = ~16'b0;
    assign data[4783] = ~16'b0;
    assign data[4784] = ~16'b0;
    assign data[4785] = ~16'b0;
    assign data[4786] = ~16'b0;
    assign data[4787] = ~16'b0;
    assign data[4788] = ~16'b0;
    assign data[4789] = ~16'b0;
    assign data[4790] = ~16'b0;
    assign data[4791] = ~16'b0;
    assign data[4792] = ~16'b0;
    assign data[4793] = ~16'b0;
    assign data[4794] = ~16'b0;
    assign data[4795] = ~16'b0;
    assign data[4796] = ~16'b0;
    assign data[4797] = ~16'b0;
    assign data[4798] = ~16'b0;
    assign data[4799] = ~16'b0;
    assign data[4800] = 16'b0;
    assign data[4801] = 16'b0;
    assign data[4802] = 16'b0;
    assign data[4803] = 16'b0;
    assign data[4804] = 16'b0;
    assign data[4805] = 16'b0;
    assign data[4806] = 16'b0;
    assign data[4807] = 16'b0;
    assign data[4808] = 16'b0;
    assign data[4809] = 16'b0;
    assign data[4810] = 16'b0;
    assign data[4811] = 16'b0;
    assign data[4812] = 16'b0;
    assign data[4813] = 16'b0;
    assign data[4814] = 16'b0;
    assign data[4815] = 16'b0;
    assign data[4816] = 16'b0;
    assign data[4817] = 16'b0;
    assign data[4818] = 16'b0;
    assign data[4819] = 16'b0;
    assign data[4820] = 16'b0;
    assign data[4821] = 16'b0;
    assign data[4822] = ~16'b0;
    assign data[4823] = ~16'b0;
    assign data[4824] = ~16'b0;
    assign data[4825] = ~16'b0;
    assign data[4826] = ~16'b0;
    assign data[4827] = ~16'b0;
    assign data[4828] = ~16'b0;
    assign data[4829] = ~16'b0;
    assign data[4830] = 16'b0;
    assign data[4831] = 16'b0;
    assign data[4832] = ~16'b0;
    assign data[4833] = ~16'b0;
    assign data[4834] = ~16'b0;
    assign data[4835] = ~16'b0;
    assign data[4836] = ~16'b0;
    assign data[4837] = ~16'b0;
    assign data[4838] = ~16'b0;
    assign data[4839] = ~16'b0;
    assign data[4840] = 16'b0;
    assign data[4841] = 16'b0;
    assign data[4842] = ~16'b0;
    assign data[4843] = ~16'b0;
    assign data[4844] = ~16'b0;
    assign data[4845] = ~16'b0;
    assign data[4846] = ~16'b0;
    assign data[4847] = ~16'b0;
    assign data[4848] = ~16'b0;
    assign data[4849] = ~16'b0;
    assign data[4850] = 16'b0;
    assign data[4851] = 16'b0;
    assign data[4852] = ~16'b0;
    assign data[4853] = ~16'b0;
    assign data[4854] = ~16'b0;
    assign data[4855] = ~16'b0;
    assign data[4856] = ~16'b0;
    assign data[4857] = ~16'b0;
    assign data[4858] = ~16'b0;
    assign data[4859] = ~16'b0;
    assign data[4860] = 16'b0;
    assign data[4861] = 16'b0;
    assign data[4862] = ~16'b0;
    assign data[4863] = ~16'b0;
    assign data[4864] = ~16'b0;
    assign data[4865] = ~16'b0;
    assign data[4866] = ~16'b0;
    assign data[4867] = ~16'b0;
    assign data[4868] = ~16'b0;
    assign data[4869] = ~16'b0;
    assign data[4870] = 16'b0;
    assign data[4871] = 16'b0;
    assign data[4872] = ~16'b0;
    assign data[4873] = ~16'b0;
    assign data[4874] = ~16'b0;
    assign data[4875] = ~16'b0;
    assign data[4876] = ~16'b0;
    assign data[4877] = ~16'b0;
    assign data[4878] = ~16'b0;
    assign data[4879] = ~16'b0;
    assign data[4880] = 16'b0;
    assign data[4881] = 16'b0;
    assign data[4882] = ~16'b0;
    assign data[4883] = ~16'b0;
    assign data[4884] = ~16'b0;
    assign data[4885] = ~16'b0;
    assign data[4886] = ~16'b0;
    assign data[4887] = ~16'b0;
    assign data[4888] = ~16'b0;
    assign data[4889] = ~16'b0;
    assign data[4890] = 16'b0;
    assign data[4891] = 16'b0;
    assign data[4892] = ~16'b0;
    assign data[4893] = ~16'b0;
    assign data[4894] = ~16'b0;
    assign data[4895] = ~16'b0;
    assign data[4896] = ~16'b0;
    assign data[4897] = ~16'b0;
    assign data[4898] = ~16'b0;
    assign data[4899] = ~16'b0;
    assign data[4900] = 16'b0;
    assign data[4901] = 16'b0;
    assign data[4902] = ~16'b0;
    assign data[4903] = ~16'b0;
    assign data[4904] = ~16'b0;
    assign data[4905] = ~16'b0;
    assign data[4906] = ~16'b0;
    assign data[4907] = ~16'b0;
    assign data[4908] = ~16'b0;
    assign data[4909] = ~16'b0;
    assign data[4910] = 16'b0;
    assign data[4911] = 16'b0;
    assign data[4912] = ~16'b0;
    assign data[4913] = ~16'b0;
    assign data[4914] = ~16'b0;
    assign data[4915] = ~16'b0;
    assign data[4916] = ~16'b0;
    assign data[4917] = ~16'b0;
    assign data[4918] = ~16'b0;
    assign data[4919] = ~16'b0;
    assign data[4920] = 16'b0;
    assign data[4921] = 16'b0;
    assign data[4922] = ~16'b0;
    assign data[4923] = ~16'b0;
    assign data[4924] = ~16'b0;
    assign data[4925] = ~16'b0;
    assign data[4926] = ~16'b0;
    assign data[4927] = ~16'b0;
    assign data[4928] = ~16'b0;
    assign data[4929] = ~16'b0;
    assign data[4930] = 16'b0;
    assign data[4931] = 16'b0;
    assign data[4932] = ~16'b0;
    assign data[4933] = ~16'b0;
    assign data[4934] = ~16'b0;
    assign data[4935] = ~16'b0;
    assign data[4936] = ~16'b0;
    assign data[4937] = ~16'b0;
    assign data[4938] = ~16'b0;
    assign data[4939] = ~16'b0;
    assign data[4940] = 16'b0;
    assign data[4941] = 16'b0;
    assign data[4942] = ~16'b0;
    assign data[4943] = ~16'b0;
    assign data[4944] = ~16'b0;
    assign data[4945] = ~16'b0;
    assign data[4946] = ~16'b0;
    assign data[4947] = ~16'b0;
    assign data[4948] = ~16'b0;
    assign data[4949] = ~16'b0;
    assign data[4950] = 16'b0;
    assign data[4951] = 16'b0;
    assign data[4952] = ~16'b0;
    assign data[4953] = ~16'b0;
    assign data[4954] = ~16'b0;
    assign data[4955] = ~16'b0;
    assign data[4956] = ~16'b0;
    assign data[4957] = ~16'b0;
    assign data[4958] = ~16'b0;
    assign data[4959] = ~16'b0;
    assign data[4960] = 16'b0;
    assign data[4961] = 16'b0;
    assign data[4962] = ~16'b0;
    assign data[4963] = ~16'b0;
    assign data[4964] = ~16'b0;
    assign data[4965] = ~16'b0;
    assign data[4966] = ~16'b0;
    assign data[4967] = ~16'b0;
    assign data[4968] = ~16'b0;
    assign data[4969] = ~16'b0;
    assign data[4970] = 16'b0;
    assign data[4971] = 16'b0;
    assign data[4972] = ~16'b0;
    assign data[4973] = ~16'b0;
    assign data[4974] = ~16'b0;
    assign data[4975] = ~16'b0;
    assign data[4976] = ~16'b0;
    assign data[4977] = ~16'b0;
    assign data[4978] = ~16'b0;
    assign data[4979] = ~16'b0;
    assign data[4980] = 16'b0;
    assign data[4981] = 16'b0;
    assign data[4982] = ~16'b0;
    assign data[4983] = ~16'b0;
    assign data[4984] = ~16'b0;
    assign data[4985] = ~16'b0;
    assign data[4986] = ~16'b0;
    assign data[4987] = ~16'b0;
    assign data[4988] = ~16'b0;
    assign data[4989] = ~16'b0;
    assign data[4990] = 16'b0;
    assign data[4991] = 16'b0;
    assign data[4992] = ~16'b0;
    assign data[4993] = ~16'b0;
    assign data[4994] = ~16'b0;
    assign data[4995] = ~16'b0;
    assign data[4996] = ~16'b0;
    assign data[4997] = ~16'b0;
    assign data[4998] = ~16'b0;
    assign data[4999] = ~16'b0;
    assign data[5000] = 16'b0;
    assign data[5001] = 16'b0;
    assign data[5002] = ~16'b0;
    assign data[5003] = ~16'b0;
    assign data[5004] = ~16'b0;
    assign data[5005] = ~16'b0;
    assign data[5006] = ~16'b0;
    assign data[5007] = ~16'b0;
    assign data[5008] = ~16'b0;
    assign data[5009] = ~16'b0;
    assign data[5010] = 16'b0;
    assign data[5011] = 16'b0;
    assign data[5012] = ~16'b0;
    assign data[5013] = ~16'b0;
    assign data[5014] = ~16'b0;
    assign data[5015] = ~16'b0;
    assign data[5016] = ~16'b0;
    assign data[5017] = ~16'b0;
    assign data[5018] = ~16'b0;
    assign data[5019] = ~16'b0;
    assign data[5020] = 16'b0;
    assign data[5021] = 16'b0;
    assign data[5022] = ~16'b0;
    assign data[5023] = ~16'b0;
    assign data[5024] = ~16'b0;
    assign data[5025] = ~16'b0;
    assign data[5026] = ~16'b0;
    assign data[5027] = ~16'b0;
    assign data[5028] = ~16'b0;
    assign data[5029] = ~16'b0;
    assign data[5030] = 16'b0;
    assign data[5031] = 16'b0;
    assign data[5032] = ~16'b0;
    assign data[5033] = ~16'b0;
    assign data[5034] = ~16'b0;
    assign data[5035] = ~16'b0;
    assign data[5036] = ~16'b0;
    assign data[5037] = ~16'b0;
    assign data[5038] = ~16'b0;
    assign data[5039] = ~16'b0;
    assign data[5040] = 16'b0;
    assign data[5041] = 16'b0;
    assign data[5042] = 16'b0;
    assign data[5043] = 16'b0;
    assign data[5044] = 16'b0;
    assign data[5045] = 16'b0;
    assign data[5046] = 16'b0;
    assign data[5047] = 16'b0;
    assign data[5048] = 16'b0;
    assign data[5049] = 16'b0;
    assign data[5050] = 16'b0;
    assign data[5051] = 16'b0;
    assign data[5052] = 16'b0;
    assign data[5053] = 16'b0;
    assign data[5054] = 16'b0;
    assign data[5055] = 16'b0;
    assign data[5056] = 16'b0;
    assign data[5057] = 16'b0;
    assign data[5058] = 16'b0;
    assign data[5059] = 16'b0;
    assign data[5060] = ~16'b0;
    assign data[5061] = ~16'b0;
    assign data[5062] = ~16'b0;
    assign data[5063] = ~16'b0;
    assign data[5064] = ~16'b0;
    assign data[5065] = ~16'b0;
    assign data[5066] = ~16'b0;
    assign data[5067] = ~16'b0;
    assign data[5068] = ~16'b0;
    assign data[5069] = ~16'b0;
    assign data[5070] = ~16'b0;
    assign data[5071] = ~16'b0;
    assign data[5072] = ~16'b0;
    assign data[5073] = ~16'b0;
    assign data[5074] = ~16'b0;
    assign data[5075] = ~16'b0;
    assign data[5076] = ~16'b0;
    assign data[5077] = ~16'b0;
    assign data[5078] = ~16'b0;
    assign data[5079] = ~16'b0;
    assign data[5080] = ~16'b0;
    assign data[5081] = ~16'b0;
    assign data[5082] = ~16'b0;
    assign data[5083] = ~16'b0;
    assign data[5084] = ~16'b0;
    assign data[5085] = ~16'b0;
    assign data[5086] = ~16'b0;
    assign data[5087] = ~16'b0;
    assign data[5088] = ~16'b0;
    assign data[5089] = ~16'b0;
    assign data[5090] = ~16'b0;
    assign data[5091] = ~16'b0;
    assign data[5092] = ~16'b0;
    assign data[5093] = ~16'b0;
    assign data[5094] = ~16'b0;
    assign data[5095] = ~16'b0;
    assign data[5096] = ~16'b0;
    assign data[5097] = ~16'b0;
    assign data[5098] = ~16'b0;
    assign data[5099] = ~16'b0;
    assign data[5100] = ~16'b0;
    assign data[5101] = ~16'b0;
    assign data[5102] = ~16'b0;
    assign data[5103] = ~16'b0;
    assign data[5104] = ~16'b0;
    assign data[5105] = ~16'b0;
    assign data[5106] = ~16'b0;
    assign data[5107] = ~16'b0;
    assign data[5108] = ~16'b0;
    assign data[5109] = ~16'b0;
    assign data[5110] = ~16'b0;
    assign data[5111] = ~16'b0;
    assign data[5112] = ~16'b0;
    assign data[5113] = ~16'b0;
    assign data[5114] = ~16'b0;
    assign data[5115] = ~16'b0;
    assign data[5116] = ~16'b0;
    assign data[5117] = ~16'b0;
    assign data[5118] = ~16'b0;
    assign data[5119] = ~16'b0;
    assign data[5120] = ~16'b0;
    assign data[5121] = ~16'b0;
    assign data[5122] = ~16'b0;
    assign data[5123] = ~16'b0;
    assign data[5124] = ~16'b0;
    assign data[5125] = ~16'b0;
    assign data[5126] = ~16'b0;
    assign data[5127] = ~16'b0;
    assign data[5128] = ~16'b0;
    assign data[5129] = ~16'b0;
    assign data[5130] = ~16'b0;
    assign data[5131] = ~16'b0;
    assign data[5132] = ~16'b0;
    assign data[5133] = ~16'b0;
    assign data[5134] = ~16'b0;
    assign data[5135] = ~16'b0;
    assign data[5136] = ~16'b0;
    assign data[5137] = ~16'b0;
    assign data[5138] = ~16'b0;
    assign data[5139] = ~16'b0;
    assign data[5140] = ~16'b0;
    assign data[5141] = ~16'b0;
    assign data[5142] = ~16'b0;
    assign data[5143] = ~16'b0;
    assign data[5144] = ~16'b0;
    assign data[5145] = ~16'b0;
    assign data[5146] = ~16'b0;
    assign data[5147] = ~16'b0;
    assign data[5148] = ~16'b0;
    assign data[5149] = ~16'b0;
    assign data[5150] = ~16'b0;
    assign data[5151] = ~16'b0;
    assign data[5152] = ~16'b0;
    assign data[5153] = ~16'b0;
    assign data[5154] = ~16'b0;
    assign data[5155] = ~16'b0;
    assign data[5156] = ~16'b0;
    assign data[5157] = ~16'b0;
    assign data[5158] = ~16'b0;
    assign data[5159] = ~16'b0;
    assign data[5160] = ~16'b0;
    assign data[5161] = ~16'b0;
    assign data[5162] = ~16'b0;
    assign data[5163] = ~16'b0;
    assign data[5164] = ~16'b0;
    assign data[5165] = ~16'b0;
    assign data[5166] = ~16'b0;
    assign data[5167] = ~16'b0;
    assign data[5168] = ~16'b0;
    assign data[5169] = ~16'b0;
    assign data[5170] = ~16'b0;
    assign data[5171] = ~16'b0;
    assign data[5172] = ~16'b0;
    assign data[5173] = ~16'b0;
    assign data[5174] = ~16'b0;
    assign data[5175] = ~16'b0;
    assign data[5176] = ~16'b0;
    assign data[5177] = ~16'b0;
    assign data[5178] = ~16'b0;
    assign data[5179] = ~16'b0;
    assign data[5180] = ~16'b0;
    assign data[5181] = ~16'b0;
    assign data[5182] = ~16'b0;
    assign data[5183] = ~16'b0;
    assign data[5184] = ~16'b0;
    assign data[5185] = ~16'b0;
    assign data[5186] = ~16'b0;
    assign data[5187] = ~16'b0;
    assign data[5188] = ~16'b0;
    assign data[5189] = ~16'b0;
    assign data[5190] = ~16'b0;
    assign data[5191] = ~16'b0;
    assign data[5192] = ~16'b0;
    assign data[5193] = ~16'b0;
    assign data[5194] = ~16'b0;
    assign data[5195] = ~16'b0;
    assign data[5196] = ~16'b0;
    assign data[5197] = ~16'b0;
    assign data[5198] = ~16'b0;
    assign data[5199] = ~16'b0;
    assign data[5200] = ~16'b0;
    assign data[5201] = ~16'b0;
    assign data[5202] = ~16'b0;
    assign data[5203] = ~16'b0;
    assign data[5204] = ~16'b0;
    assign data[5205] = ~16'b0;
    assign data[5206] = ~16'b0;
    assign data[5207] = ~16'b0;
    assign data[5208] = ~16'b0;
    assign data[5209] = ~16'b0;
    assign data[5210] = ~16'b0;
    assign data[5211] = ~16'b0;
    assign data[5212] = ~16'b0;
    assign data[5213] = ~16'b0;
    assign data[5214] = ~16'b0;
    assign data[5215] = ~16'b0;
    assign data[5216] = ~16'b0;
    assign data[5217] = ~16'b0;
    assign data[5218] = ~16'b0;
    assign data[5219] = ~16'b0;
    assign data[5220] = ~16'b0;
    assign data[5221] = ~16'b0;
    assign data[5222] = ~16'b0;
    assign data[5223] = ~16'b0;
    assign data[5224] = ~16'b0;
    assign data[5225] = ~16'b0;
    assign data[5226] = ~16'b0;
    assign data[5227] = ~16'b0;
    assign data[5228] = ~16'b0;
    assign data[5229] = ~16'b0;
    assign data[5230] = 16'b0;
    assign data[5231] = 16'b0;
    assign data[5232] = 16'b0;
    assign data[5233] = 16'b0;
    assign data[5234] = 16'b0;
    assign data[5235] = 16'b0;
    assign data[5236] = 16'b0;
    assign data[5237] = 16'b0;
    assign data[5238] = 16'b0;
    assign data[5239] = 16'b0;
    assign data[5240] = 16'b0;
    assign data[5241] = 16'b0;
    assign data[5242] = 16'b0;
    assign data[5243] = 16'b0;
    assign data[5244] = 16'b0;
    assign data[5245] = 16'b0;
    assign data[5246] = 16'b0;
    assign data[5247] = 16'b0;
    assign data[5248] = 16'b0;
    assign data[5249] = 16'b0;
    assign data[5250] = 16'b0;
    assign data[5251] = 16'b0;
    assign data[5252] = ~16'b0;
    assign data[5253] = ~16'b0;
    assign data[5254] = ~16'b0;
    assign data[5255] = ~16'b0;
    assign data[5256] = ~16'b0;
    assign data[5257] = ~16'b0;
    assign data[5258] = ~16'b0;
    assign data[5259] = ~16'b0;
    assign data[5260] = 16'b0;
    assign data[5261] = 16'b0;
    assign data[5262] = ~16'b0;
    assign data[5263] = ~16'b0;
    assign data[5264] = ~16'b0;
    assign data[5265] = ~16'b0;
    assign data[5266] = ~16'b0;
    assign data[5267] = ~16'b0;
    assign data[5268] = ~16'b0;
    assign data[5269] = ~16'b0;
    assign data[5270] = 16'b0;
    assign data[5271] = 16'b0;
    assign data[5272] = ~16'b0;
    assign data[5273] = ~16'b0;
    assign data[5274] = ~16'b0;
    assign data[5275] = ~16'b0;
    assign data[5276] = ~16'b0;
    assign data[5277] = ~16'b0;
    assign data[5278] = ~16'b0;
    assign data[5279] = ~16'b0;
    assign data[5280] = 16'b0;
    assign data[5281] = 16'b0;
    assign data[5282] = ~16'b0;
    assign data[5283] = ~16'b0;
    assign data[5284] = ~16'b0;
    assign data[5285] = ~16'b0;
    assign data[5286] = ~16'b0;
    assign data[5287] = ~16'b0;
    assign data[5288] = ~16'b0;
    assign data[5289] = ~16'b0;
    assign data[5290] = 16'b0;
    assign data[5291] = 16'b0;
    assign data[5292] = ~16'b0;
    assign data[5293] = ~16'b0;
    assign data[5294] = ~16'b0;
    assign data[5295] = ~16'b0;
    assign data[5296] = ~16'b0;
    assign data[5297] = ~16'b0;
    assign data[5298] = ~16'b0;
    assign data[5299] = ~16'b0;
    assign data[5300] = 16'b0;
    assign data[5301] = 16'b0;
    assign data[5302] = ~16'b0;
    assign data[5303] = ~16'b0;
    assign data[5304] = ~16'b0;
    assign data[5305] = ~16'b0;
    assign data[5306] = ~16'b0;
    assign data[5307] = ~16'b0;
    assign data[5308] = ~16'b0;
    assign data[5309] = ~16'b0;
    assign data[5310] = 16'b0;
    assign data[5311] = 16'b0;
    assign data[5312] = ~16'b0;
    assign data[5313] = ~16'b0;
    assign data[5314] = ~16'b0;
    assign data[5315] = ~16'b0;
    assign data[5316] = ~16'b0;
    assign data[5317] = ~16'b0;
    assign data[5318] = ~16'b0;
    assign data[5319] = ~16'b0;
    assign data[5320] = 16'b0;
    assign data[5321] = 16'b0;
    assign data[5322] = ~16'b0;
    assign data[5323] = ~16'b0;
    assign data[5324] = ~16'b0;
    assign data[5325] = ~16'b0;
    assign data[5326] = ~16'b0;
    assign data[5327] = ~16'b0;
    assign data[5328] = ~16'b0;
    assign data[5329] = ~16'b0;
    assign data[5330] = 16'b0;
    assign data[5331] = 16'b0;
    assign data[5332] = ~16'b0;
    assign data[5333] = ~16'b0;
    assign data[5334] = ~16'b0;
    assign data[5335] = ~16'b0;
    assign data[5336] = ~16'b0;
    assign data[5337] = ~16'b0;
    assign data[5338] = ~16'b0;
    assign data[5339] = ~16'b0;
    assign data[5340] = 16'b0;
    assign data[5341] = 16'b0;
    assign data[5342] = ~16'b0;
    assign data[5343] = ~16'b0;
    assign data[5344] = ~16'b0;
    assign data[5345] = ~16'b0;
    assign data[5346] = ~16'b0;
    assign data[5347] = ~16'b0;
    assign data[5348] = ~16'b0;
    assign data[5349] = ~16'b0;
    assign data[5350] = 16'b0;
    assign data[5351] = 16'b0;
    assign data[5352] = ~16'b0;
    assign data[5353] = ~16'b0;
    assign data[5354] = ~16'b0;
    assign data[5355] = ~16'b0;
    assign data[5356] = ~16'b0;
    assign data[5357] = ~16'b0;
    assign data[5358] = ~16'b0;
    assign data[5359] = ~16'b0;
    assign data[5360] = 16'b0;
    assign data[5361] = 16'b0;
    assign data[5362] = ~16'b0;
    assign data[5363] = ~16'b0;
    assign data[5364] = ~16'b0;
    assign data[5365] = ~16'b0;
    assign data[5366] = ~16'b0;
    assign data[5367] = ~16'b0;
    assign data[5368] = ~16'b0;
    assign data[5369] = ~16'b0;
    assign data[5370] = 16'b0;
    assign data[5371] = 16'b0;
    assign data[5372] = ~16'b0;
    assign data[5373] = ~16'b0;
    assign data[5374] = ~16'b0;
    assign data[5375] = ~16'b0;
    assign data[5376] = ~16'b0;
    assign data[5377] = ~16'b0;
    assign data[5378] = ~16'b0;
    assign data[5379] = ~16'b0;
    assign data[5380] = 16'b0;
    assign data[5381] = 16'b0;
    assign data[5382] = ~16'b0;
    assign data[5383] = ~16'b0;
    assign data[5384] = ~16'b0;
    assign data[5385] = ~16'b0;
    assign data[5386] = ~16'b0;
    assign data[5387] = ~16'b0;
    assign data[5388] = ~16'b0;
    assign data[5389] = ~16'b0;
    assign data[5390] = 16'b0;
    assign data[5391] = 16'b0;
    assign data[5392] = ~16'b0;
    assign data[5393] = ~16'b0;
    assign data[5394] = ~16'b0;
    assign data[5395] = ~16'b0;
    assign data[5396] = ~16'b0;
    assign data[5397] = ~16'b0;
    assign data[5398] = ~16'b0;
    assign data[5399] = ~16'b0;
    assign data[5400] = 16'b0;
    assign data[5401] = 16'b0;
    assign data[5402] = ~16'b0;
    assign data[5403] = ~16'b0;
    assign data[5404] = ~16'b0;
    assign data[5405] = ~16'b0;
    assign data[5406] = ~16'b0;
    assign data[5407] = ~16'b0;
    assign data[5408] = ~16'b0;
    assign data[5409] = ~16'b0;
    assign data[5410] = 16'b0;
    assign data[5411] = 16'b0;
    assign data[5412] = ~16'b0;
    assign data[5413] = ~16'b0;
    assign data[5414] = ~16'b0;
    assign data[5415] = ~16'b0;
    assign data[5416] = ~16'b0;
    assign data[5417] = ~16'b0;
    assign data[5418] = ~16'b0;
    assign data[5419] = ~16'b0;
    assign data[5420] = 16'b0;
    assign data[5421] = 16'b0;
    assign data[5422] = ~16'b0;
    assign data[5423] = ~16'b0;
    assign data[5424] = ~16'b0;
    assign data[5425] = ~16'b0;
    assign data[5426] = ~16'b0;
    assign data[5427] = ~16'b0;
    assign data[5428] = ~16'b0;
    assign data[5429] = ~16'b0;
    assign data[5430] = 16'b0;
    assign data[5431] = 16'b0;
    assign data[5432] = ~16'b0;
    assign data[5433] = ~16'b0;
    assign data[5434] = ~16'b0;
    assign data[5435] = ~16'b0;
    assign data[5436] = ~16'b0;
    assign data[5437] = ~16'b0;
    assign data[5438] = ~16'b0;
    assign data[5439] = ~16'b0;
    assign data[5440] = 16'b0;
    assign data[5441] = 16'b0;
    assign data[5442] = ~16'b0;
    assign data[5443] = ~16'b0;
    assign data[5444] = ~16'b0;
    assign data[5445] = ~16'b0;
    assign data[5446] = ~16'b0;
    assign data[5447] = ~16'b0;
    assign data[5448] = ~16'b0;
    assign data[5449] = ~16'b0;
    assign data[5450] = 16'b0;
    assign data[5451] = 16'b0;
    assign data[5452] = ~16'b0;
    assign data[5453] = ~16'b0;
    assign data[5454] = ~16'b0;
    assign data[5455] = ~16'b0;
    assign data[5456] = ~16'b0;
    assign data[5457] = ~16'b0;
    assign data[5458] = ~16'b0;
    assign data[5459] = ~16'b0;
    assign data[5460] = 16'b0;
    assign data[5461] = 16'b0;
    assign data[5462] = ~16'b0;
    assign data[5463] = ~16'b0;
    assign data[5464] = ~16'b0;
    assign data[5465] = ~16'b0;
    assign data[5466] = ~16'b0;
    assign data[5467] = ~16'b0;
    assign data[5468] = ~16'b0;
    assign data[5469] = ~16'b0;
    assign data[5470] = 16'b0;
    assign data[5471] = 16'b0;
    assign data[5472] = ~16'b0;
    assign data[5473] = ~16'b0;
    assign data[5474] = ~16'b0;
    assign data[5475] = ~16'b0;
    assign data[5476] = ~16'b0;
    assign data[5477] = ~16'b0;
    assign data[5478] = ~16'b0;
    assign data[5479] = ~16'b0;
    assign data[5480] = 16'b0;
    assign data[5481] = 16'b0;
    assign data[5482] = ~16'b0;
    assign data[5483] = ~16'b0;
    assign data[5484] = ~16'b0;
    assign data[5485] = ~16'b0;
    assign data[5486] = ~16'b0;
    assign data[5487] = ~16'b0;
    assign data[5488] = ~16'b0;
    assign data[5489] = ~16'b0;
    assign data[5490] = 16'b0;
    assign data[5491] = 16'b0;
    assign data[5492] = ~16'b0;
    assign data[5493] = ~16'b0;
    assign data[5494] = ~16'b0;
    assign data[5495] = ~16'b0;
    assign data[5496] = ~16'b0;
    assign data[5497] = ~16'b0;
    assign data[5498] = ~16'b0;
    assign data[5499] = ~16'b0;
    assign data[5500] = 16'b0;
    assign data[5501] = 16'b0;
    assign data[5502] = ~16'b0;
    assign data[5503] = ~16'b0;
    assign data[5504] = ~16'b0;
    assign data[5505] = ~16'b0;
    assign data[5506] = ~16'b0;
    assign data[5507] = ~16'b0;
    assign data[5508] = ~16'b0;
    assign data[5509] = ~16'b0;
    assign data[5510] = 16'b0;
    assign data[5511] = 16'b0;
    assign data[5512] = ~16'b0;
    assign data[5513] = ~16'b0;
    assign data[5514] = ~16'b0;
    assign data[5515] = ~16'b0;
    assign data[5516] = ~16'b0;
    assign data[5517] = ~16'b0;
    assign data[5518] = ~16'b0;
    assign data[5519] = ~16'b0;
    assign data[5520] = 16'b0;
    assign data[5521] = 16'b0;
    assign data[5522] = ~16'b0;
    assign data[5523] = ~16'b0;
    assign data[5524] = ~16'b0;
    assign data[5525] = ~16'b0;
    assign data[5526] = ~16'b0;
    assign data[5527] = ~16'b0;
    assign data[5528] = ~16'b0;
    assign data[5529] = ~16'b0;
    assign data[5530] = 16'b0;
    assign data[5531] = 16'b0;
    assign data[5532] = ~16'b0;
    assign data[5533] = ~16'b0;
    assign data[5534] = ~16'b0;
    assign data[5535] = ~16'b0;
    assign data[5536] = ~16'b0;
    assign data[5537] = ~16'b0;
    assign data[5538] = ~16'b0;
    assign data[5539] = ~16'b0;
    assign data[5540] = 16'b0;
    assign data[5541] = 16'b0;
    assign data[5542] = ~16'b0;
    assign data[5543] = ~16'b0;
    assign data[5544] = ~16'b0;
    assign data[5545] = ~16'b0;
    assign data[5546] = ~16'b0;
    assign data[5547] = ~16'b0;
    assign data[5548] = ~16'b0;
    assign data[5549] = ~16'b0;
    assign data[5550] = 16'b0;
    assign data[5551] = 16'b0;
    assign data[5552] = ~16'b0;
    assign data[5553] = ~16'b0;
    assign data[5554] = ~16'b0;
    assign data[5555] = ~16'b0;
    assign data[5556] = ~16'b0;
    assign data[5557] = ~16'b0;
    assign data[5558] = ~16'b0;
    assign data[5559] = ~16'b0;
    assign data[5560] = 16'b0;
    assign data[5561] = 16'b0;
    assign data[5562] = ~16'b0;
    assign data[5563] = ~16'b0;
    assign data[5564] = ~16'b0;
    assign data[5565] = ~16'b0;
    assign data[5566] = ~16'b0;
    assign data[5567] = ~16'b0;
    assign data[5568] = ~16'b0;
    assign data[5569] = ~16'b0;
    assign data[5570] = 16'b0;
    assign data[5571] = 16'b0;
    assign data[5572] = ~16'b0;
    assign data[5573] = ~16'b0;
    assign data[5574] = ~16'b0;
    assign data[5575] = ~16'b0;
    assign data[5576] = ~16'b0;
    assign data[5577] = ~16'b0;
    assign data[5578] = ~16'b0;
    assign data[5579] = ~16'b0;
    assign data[5580] = 16'b0;
    assign data[5581] = 16'b0;
    assign data[5582] = ~16'b0;
    assign data[5583] = ~16'b0;
    assign data[5584] = ~16'b0;
    assign data[5585] = ~16'b0;
    assign data[5586] = ~16'b0;
    assign data[5587] = ~16'b0;
    assign data[5588] = ~16'b0;
    assign data[5589] = ~16'b0;
    assign data[5590] = 16'b0;
    assign data[5591] = 16'b0;
    assign data[5592] = ~16'b0;
    assign data[5593] = ~16'b0;
    assign data[5594] = ~16'b0;
    assign data[5595] = ~16'b0;
    assign data[5596] = ~16'b0;
    assign data[5597] = ~16'b0;
    assign data[5598] = ~16'b0;
    assign data[5599] = ~16'b0;
    assign data[5600] = 16'b0;
    assign data[5601] = 16'b0;
    assign data[5602] = ~16'b0;
    assign data[5603] = ~16'b0;
    assign data[5604] = ~16'b0;
    assign data[5605] = ~16'b0;
    assign data[5606] = ~16'b0;
    assign data[5607] = ~16'b0;
    assign data[5608] = ~16'b0;
    assign data[5609] = ~16'b0;
    assign data[5610] = 16'b0;
    assign data[5611] = 16'b0;
    assign data[5612] = 16'b0;
    assign data[5613] = 16'b0;
    assign data[5614] = 16'b0;
    assign data[5615] = 16'b0;
    assign data[5616] = 16'b0;
    assign data[5617] = 16'b0;
    assign data[5618] = 16'b0;
    assign data[5619] = 16'b0;
    assign data[5620] = 16'b0;
    assign data[5621] = 16'b0;
    assign data[5622] = 16'b0;
    assign data[5623] = 16'b0;
    assign data[5624] = 16'b0;
    assign data[5625] = 16'b0;
    assign data[5626] = 16'b0;
    assign data[5627] = 16'b0;
    assign data[5628] = 16'b0;
    assign data[5629] = 16'b0;
    assign data[5630] = ~16'b0;
    assign data[5631] = ~16'b0;
    assign data[5632] = ~16'b0;
    assign data[5633] = ~16'b0;
    assign data[5634] = ~16'b0;
    assign data[5635] = ~16'b0;
    assign data[5636] = ~16'b0;
    assign data[5637] = ~16'b0;
    assign data[5638] = ~16'b0;
    assign data[5639] = ~16'b0;
    assign data[5640] = ~16'b0;
    assign data[5641] = ~16'b0;
    assign data[5642] = ~16'b0;
    assign data[5643] = ~16'b0;
    assign data[5644] = ~16'b0;
    assign data[5645] = ~16'b0;
    assign data[5646] = ~16'b0;
    assign data[5647] = ~16'b0;
    assign data[5648] = ~16'b0;
    assign data[5649] = ~16'b0;
    assign data[5650] = ~16'b0;
    assign data[5651] = ~16'b0;
    assign data[5652] = ~16'b0;
    assign data[5653] = ~16'b0;
    assign data[5654] = ~16'b0;
    assign data[5655] = ~16'b0;
    assign data[5656] = ~16'b0;
    assign data[5657] = ~16'b0;
    assign data[5658] = ~16'b0;
    assign data[5659] = ~16'b0;
    assign data[5660] = ~16'b0;
    assign data[5661] = ~16'b0;
    assign data[5662] = ~16'b0;
    assign data[5663] = ~16'b0;
    assign data[5664] = ~16'b0;
    assign data[5665] = ~16'b0;
    assign data[5666] = ~16'b0;
    assign data[5667] = ~16'b0;
    assign data[5668] = ~16'b0;
    assign data[5669] = ~16'b0;
    assign data[5670] = ~16'b0;
    assign data[5671] = ~16'b0;
    assign data[5672] = ~16'b0;
    assign data[5673] = ~16'b0;
    assign data[5674] = ~16'b0;
    assign data[5675] = ~16'b0;
    assign data[5676] = ~16'b0;
    assign data[5677] = ~16'b0;
    assign data[5678] = ~16'b0;
    assign data[5679] = ~16'b0;
    assign data[5680] = ~16'b0;
    assign data[5681] = ~16'b0;
    assign data[5682] = ~16'b0;
    assign data[5683] = ~16'b0;
    assign data[5684] = ~16'b0;
    assign data[5685] = ~16'b0;
    assign data[5686] = ~16'b0;
    assign data[5687] = ~16'b0;
    assign data[5688] = ~16'b0;
    assign data[5689] = ~16'b0;
    assign data[5690] = ~16'b0;
    assign data[5691] = ~16'b0;
    assign data[5692] = ~16'b0;
    assign data[5693] = ~16'b0;
    assign data[5694] = ~16'b0;
    assign data[5695] = ~16'b0;
    assign data[5696] = ~16'b0;
    assign data[5697] = ~16'b0;
    assign data[5698] = ~16'b0;
    assign data[5699] = ~16'b0;
    assign data[5700] = ~16'b0;
    assign data[5701] = ~16'b0;
    assign data[5702] = ~16'b0;
    assign data[5703] = ~16'b0;
    assign data[5704] = ~16'b0;
    assign data[5705] = ~16'b0;
    assign data[5706] = ~16'b0;
    assign data[5707] = ~16'b0;
    assign data[5708] = ~16'b0;
    assign data[5709] = ~16'b0;
    assign data[5710] = ~16'b0;
    assign data[5711] = ~16'b0;
    assign data[5712] = ~16'b0;
    assign data[5713] = ~16'b0;
    assign data[5714] = ~16'b0;
    assign data[5715] = ~16'b0;
    assign data[5716] = ~16'b0;
    assign data[5717] = ~16'b0;
    assign data[5718] = ~16'b0;
    assign data[5719] = ~16'b0;
    assign data[5720] = ~16'b0;
    assign data[5721] = ~16'b0;
    assign data[5722] = ~16'b0;
    assign data[5723] = ~16'b0;
    assign data[5724] = ~16'b0;
    assign data[5725] = ~16'b0;
    assign data[5726] = ~16'b0;
    assign data[5727] = ~16'b0;
    assign data[5728] = ~16'b0;
    assign data[5729] = ~16'b0;
    assign data[5730] = ~16'b0;
    assign data[5731] = ~16'b0;
    assign data[5732] = ~16'b0;
    assign data[5733] = ~16'b0;
    assign data[5734] = ~16'b0;
    assign data[5735] = ~16'b0;
    assign data[5736] = ~16'b0;
    assign data[5737] = ~16'b0;
    assign data[5738] = ~16'b0;
    assign data[5739] = ~16'b0;
    assign data[5740] = ~16'b0;
    assign data[5741] = ~16'b0;
    assign data[5742] = ~16'b0;
    assign data[5743] = ~16'b0;
    assign data[5744] = ~16'b0;
    assign data[5745] = ~16'b0;
    assign data[5746] = ~16'b0;
    assign data[5747] = ~16'b0;
    assign data[5748] = ~16'b0;
    assign data[5749] = ~16'b0;
    assign data[5750] = ~16'b0;
    assign data[5751] = ~16'b0;
    assign data[5752] = ~16'b0;
    assign data[5753] = ~16'b0;
    assign data[5754] = ~16'b0;
    assign data[5755] = ~16'b0;
    assign data[5756] = ~16'b0;
    assign data[5757] = ~16'b0;
    assign data[5758] = ~16'b0;
    assign data[5759] = ~16'b0;
    assign data[5760] = ~16'b0;
    assign data[5761] = ~16'b0;
    assign data[5762] = ~16'b0;
    assign data[5763] = ~16'b0;
    assign data[5764] = ~16'b0;
    assign data[5765] = ~16'b0;
    assign data[5766] = ~16'b0;
    assign data[5767] = ~16'b0;
    assign data[5768] = ~16'b0;
    assign data[5769] = ~16'b0;
    assign data[5770] = ~16'b0;
    assign data[5771] = ~16'b0;
    assign data[5772] = ~16'b0;
    assign data[5773] = ~16'b0;
    assign data[5774] = ~16'b0;
    assign data[5775] = ~16'b0;
    assign data[5776] = ~16'b0;
    assign data[5777] = ~16'b0;
    assign data[5778] = ~16'b0;
    assign data[5779] = ~16'b0;
    assign data[5780] = ~16'b0;
    assign data[5781] = ~16'b0;
    assign data[5782] = ~16'b0;
    assign data[5783] = ~16'b0;
    assign data[5784] = ~16'b0;
    assign data[5785] = ~16'b0;
    assign data[5786] = ~16'b0;
    assign data[5787] = ~16'b0;
    assign data[5788] = ~16'b0;
    assign data[5789] = ~16'b0;
    assign data[5790] = ~16'b0;
    assign data[5791] = ~16'b0;
    assign data[5792] = ~16'b0;
    assign data[5793] = ~16'b0;
    assign data[5794] = ~16'b0;
    assign data[5795] = ~16'b0;
    assign data[5796] = ~16'b0;
    assign data[5797] = ~16'b0;
    assign data[5798] = ~16'b0;
    assign data[5799] = ~16'b0;
    assign data[5800] = 16'b0;
    assign data[5801] = 16'b0;
    assign data[5802] = 16'b0;
    assign data[5803] = 16'b0;
    assign data[5804] = 16'b0;
    assign data[5805] = 16'b0;
    assign data[5806] = 16'b0;
    assign data[5807] = 16'b0;
    assign data[5808] = 16'b0;
    assign data[5809] = 16'b0;
    assign data[5810] = 16'b0;
    assign data[5811] = 16'b0;
    assign data[5812] = 16'b0;
    assign data[5813] = 16'b0;
    assign data[5814] = 16'b0;
    assign data[5815] = 16'b0;
    assign data[5816] = 16'b0;
    assign data[5817] = 16'b0;
    assign data[5818] = 16'b0;
    assign data[5819] = 16'b0;
    assign data[5820] = 16'b0;
    assign data[5821] = 16'b0;
    assign data[5822] = ~16'b0;
    assign data[5823] = ~16'b0;
    assign data[5824] = ~16'b0;
    assign data[5825] = ~16'b0;
    assign data[5826] = ~16'b0;
    assign data[5827] = ~16'b0;
    assign data[5828] = ~16'b0;
    assign data[5829] = ~16'b0;
    assign data[5830] = 16'b0;
    assign data[5831] = 16'b0;
    assign data[5832] = ~16'b0;
    assign data[5833] = ~16'b0;
    assign data[5834] = ~16'b0;
    assign data[5835] = ~16'b0;
    assign data[5836] = ~16'b0;
    assign data[5837] = ~16'b0;
    assign data[5838] = ~16'b0;
    assign data[5839] = ~16'b0;
    assign data[5840] = 16'b0;
    assign data[5841] = 16'b0;
    assign data[5842] = ~16'b0;
    assign data[5843] = ~16'b0;
    assign data[5844] = ~16'b0;
    assign data[5845] = ~16'b0;
    assign data[5846] = ~16'b0;
    assign data[5847] = ~16'b0;
    assign data[5848] = ~16'b0;
    assign data[5849] = ~16'b0;
    assign data[5850] = 16'b0;
    assign data[5851] = 16'b0;
    assign data[5852] = ~16'b0;
    assign data[5853] = ~16'b0;
    assign data[5854] = ~16'b0;
    assign data[5855] = ~16'b0;
    assign data[5856] = ~16'b0;
    assign data[5857] = ~16'b0;
    assign data[5858] = ~16'b0;
    assign data[5859] = ~16'b0;
    assign data[5860] = 16'b0;
    assign data[5861] = 16'b0;
    assign data[5862] = ~16'b0;
    assign data[5863] = ~16'b0;
    assign data[5864] = ~16'b0;
    assign data[5865] = ~16'b0;
    assign data[5866] = ~16'b0;
    assign data[5867] = ~16'b0;
    assign data[5868] = ~16'b0;
    assign data[5869] = ~16'b0;
    assign data[5870] = 16'b0;
    assign data[5871] = 16'b0;
    assign data[5872] = ~16'b0;
    assign data[5873] = ~16'b0;
    assign data[5874] = ~16'b0;
    assign data[5875] = ~16'b0;
    assign data[5876] = ~16'b0;
    assign data[5877] = ~16'b0;
    assign data[5878] = ~16'b0;
    assign data[5879] = ~16'b0;
    assign data[5880] = 16'b0;
    assign data[5881] = 16'b0;
    assign data[5882] = ~16'b0;
    assign data[5883] = ~16'b0;
    assign data[5884] = ~16'b0;
    assign data[5885] = ~16'b0;
    assign data[5886] = ~16'b0;
    assign data[5887] = ~16'b0;
    assign data[5888] = ~16'b0;
    assign data[5889] = ~16'b0;
    assign data[5890] = 16'b0;
    assign data[5891] = 16'b0;
    assign data[5892] = ~16'b0;
    assign data[5893] = ~16'b0;
    assign data[5894] = ~16'b0;
    assign data[5895] = ~16'b0;
    assign data[5896] = ~16'b0;
    assign data[5897] = ~16'b0;
    assign data[5898] = ~16'b0;
    assign data[5899] = ~16'b0;
    assign data[5900] = 16'b0;
    assign data[5901] = 16'b0;
    assign data[5902] = ~16'b0;
    assign data[5903] = ~16'b0;
    assign data[5904] = ~16'b0;
    assign data[5905] = ~16'b0;
    assign data[5906] = ~16'b0;
    assign data[5907] = ~16'b0;
    assign data[5908] = ~16'b0;
    assign data[5909] = ~16'b0;
    assign data[5910] = 16'b0;
    assign data[5911] = 16'b0;
    assign data[5912] = ~16'b0;
    assign data[5913] = ~16'b0;
    assign data[5914] = ~16'b0;
    assign data[5915] = ~16'b0;
    assign data[5916] = ~16'b0;
    assign data[5917] = ~16'b0;
    assign data[5918] = ~16'b0;
    assign data[5919] = ~16'b0;
    assign data[5920] = 16'b0;
    assign data[5921] = 16'b0;
    assign data[5922] = ~16'b0;
    assign data[5923] = ~16'b0;
    assign data[5924] = ~16'b0;
    assign data[5925] = ~16'b0;
    assign data[5926] = ~16'b0;
    assign data[5927] = ~16'b0;
    assign data[5928] = ~16'b0;
    assign data[5929] = ~16'b0;
    assign data[5930] = 16'b0;
    assign data[5931] = 16'b0;
    assign data[5932] = ~16'b0;
    assign data[5933] = ~16'b0;
    assign data[5934] = ~16'b0;
    assign data[5935] = ~16'b0;
    assign data[5936] = ~16'b0;
    assign data[5937] = ~16'b0;
    assign data[5938] = ~16'b0;
    assign data[5939] = ~16'b0;
    assign data[5940] = 16'b0;
    assign data[5941] = 16'b0;
    assign data[5942] = ~16'b0;
    assign data[5943] = ~16'b0;
    assign data[5944] = ~16'b0;
    assign data[5945] = ~16'b0;
    assign data[5946] = ~16'b0;
    assign data[5947] = ~16'b0;
    assign data[5948] = ~16'b0;
    assign data[5949] = ~16'b0;
    assign data[5950] = 16'b0;
    assign data[5951] = 16'b0;
    assign data[5952] = ~16'b0;
    assign data[5953] = ~16'b0;
    assign data[5954] = ~16'b0;
    assign data[5955] = ~16'b0;
    assign data[5956] = ~16'b0;
    assign data[5957] = ~16'b0;
    assign data[5958] = ~16'b0;
    assign data[5959] = ~16'b0;
    assign data[5960] = 16'b0;
    assign data[5961] = 16'b0;
    assign data[5962] = ~16'b0;
    assign data[5963] = ~16'b0;
    assign data[5964] = ~16'b0;
    assign data[5965] = ~16'b0;
    assign data[5966] = ~16'b0;
    assign data[5967] = ~16'b0;
    assign data[5968] = ~16'b0;
    assign data[5969] = ~16'b0;
    assign data[5970] = 16'b0;
    assign data[5971] = 16'b0;
    assign data[5972] = ~16'b0;
    assign data[5973] = ~16'b0;
    assign data[5974] = ~16'b0;
    assign data[5975] = ~16'b0;
    assign data[5976] = ~16'b0;
    assign data[5977] = ~16'b0;
    assign data[5978] = ~16'b0;
    assign data[5979] = ~16'b0;
    assign data[5980] = 16'b0;
    assign data[5981] = 16'b0;
    assign data[5982] = ~16'b0;
    assign data[5983] = ~16'b0;
    assign data[5984] = ~16'b0;
    assign data[5985] = ~16'b0;
    assign data[5986] = ~16'b0;
    assign data[5987] = ~16'b0;
    assign data[5988] = ~16'b0;
    assign data[5989] = ~16'b0;
    assign data[5990] = 16'b0;
    assign data[5991] = 16'b0;
    assign data[5992] = ~16'b0;
    assign data[5993] = ~16'b0;
    assign data[5994] = ~16'b0;
    assign data[5995] = ~16'b0;
    assign data[5996] = ~16'b0;
    assign data[5997] = ~16'b0;
    assign data[5998] = ~16'b0;
    assign data[5999] = ~16'b0;
    assign data[6000] = 16'b0;
    assign data[6001] = 16'b0;
    assign data[6002] = ~16'b0;
    assign data[6003] = ~16'b0;
    assign data[6004] = ~16'b0;
    assign data[6005] = ~16'b0;
    assign data[6006] = ~16'b0;
    assign data[6007] = ~16'b0;
    assign data[6008] = ~16'b0;
    assign data[6009] = ~16'b0;
    assign data[6010] = 16'b0;
    assign data[6011] = 16'b0;
    assign data[6012] = ~16'b0;
    assign data[6013] = ~16'b0;
    assign data[6014] = ~16'b0;
    assign data[6015] = ~16'b0;
    assign data[6016] = ~16'b0;
    assign data[6017] = ~16'b0;
    assign data[6018] = ~16'b0;
    assign data[6019] = ~16'b0;
    assign data[6020] = 16'b0;
    assign data[6021] = 16'b0;
    assign data[6022] = ~16'b0;
    assign data[6023] = ~16'b0;
    assign data[6024] = ~16'b0;
    assign data[6025] = ~16'b0;
    assign data[6026] = ~16'b0;
    assign data[6027] = ~16'b0;
    assign data[6028] = ~16'b0;
    assign data[6029] = ~16'b0;
    assign data[6030] = 16'b0;
    assign data[6031] = 16'b0;
    assign data[6032] = ~16'b0;
    assign data[6033] = ~16'b0;
    assign data[6034] = ~16'b0;
    assign data[6035] = ~16'b0;
    assign data[6036] = ~16'b0;
    assign data[6037] = ~16'b0;
    assign data[6038] = ~16'b0;
    assign data[6039] = ~16'b0;
    assign data[6040] = 16'b0;
    assign data[6041] = 16'b0;
    assign data[6042] = ~16'b0;
    assign data[6043] = ~16'b0;
    assign data[6044] = ~16'b0;
    assign data[6045] = ~16'b0;
    assign data[6046] = ~16'b0;
    assign data[6047] = ~16'b0;
    assign data[6048] = ~16'b0;
    assign data[6049] = ~16'b0;
    assign data[6050] = 16'b0;
    assign data[6051] = 16'b0;
    assign data[6052] = ~16'b0;
    assign data[6053] = ~16'b0;
    assign data[6054] = ~16'b0;
    assign data[6055] = ~16'b0;
    assign data[6056] = ~16'b0;
    assign data[6057] = ~16'b0;
    assign data[6058] = ~16'b0;
    assign data[6059] = ~16'b0;
    assign data[6060] = 16'b0;
    assign data[6061] = 16'b0;
    assign data[6062] = ~16'b0;
    assign data[6063] = ~16'b0;
    assign data[6064] = ~16'b0;
    assign data[6065] = ~16'b0;
    assign data[6066] = ~16'b0;
    assign data[6067] = ~16'b0;
    assign data[6068] = ~16'b0;
    assign data[6069] = ~16'b0;
    assign data[6070] = 16'b0;
    assign data[6071] = 16'b0;
    assign data[6072] = ~16'b0;
    assign data[6073] = ~16'b0;
    assign data[6074] = ~16'b0;
    assign data[6075] = ~16'b0;
    assign data[6076] = ~16'b0;
    assign data[6077] = ~16'b0;
    assign data[6078] = ~16'b0;
    assign data[6079] = ~16'b0;
    assign data[6080] = 16'b0;
    assign data[6081] = 16'b0;
    assign data[6082] = ~16'b0;
    assign data[6083] = ~16'b0;
    assign data[6084] = ~16'b0;
    assign data[6085] = ~16'b0;
    assign data[6086] = ~16'b0;
    assign data[6087] = ~16'b0;
    assign data[6088] = ~16'b0;
    assign data[6089] = ~16'b0;
    assign data[6090] = 16'b0;
    assign data[6091] = 16'b0;
    assign data[6092] = ~16'b0;
    assign data[6093] = ~16'b0;
    assign data[6094] = ~16'b0;
    assign data[6095] = ~16'b0;
    assign data[6096] = ~16'b0;
    assign data[6097] = ~16'b0;
    assign data[6098] = ~16'b0;
    assign data[6099] = ~16'b0;
    assign data[6100] = 16'b0;
    assign data[6101] = 16'b0;
    assign data[6102] = ~16'b0;
    assign data[6103] = ~16'b0;
    assign data[6104] = ~16'b0;
    assign data[6105] = ~16'b0;
    assign data[6106] = ~16'b0;
    assign data[6107] = ~16'b0;
    assign data[6108] = ~16'b0;
    assign data[6109] = ~16'b0;
    assign data[6110] = 16'b0;
    assign data[6111] = 16'b0;
    assign data[6112] = ~16'b0;
    assign data[6113] = ~16'b0;
    assign data[6114] = ~16'b0;
    assign data[6115] = ~16'b0;
    assign data[6116] = ~16'b0;
    assign data[6117] = ~16'b0;
    assign data[6118] = ~16'b0;
    assign data[6119] = ~16'b0;
    assign data[6120] = 16'b0;
    assign data[6121] = 16'b0;
    assign data[6122] = ~16'b0;
    assign data[6123] = ~16'b0;
    assign data[6124] = ~16'b0;
    assign data[6125] = ~16'b0;
    assign data[6126] = ~16'b0;
    assign data[6127] = ~16'b0;
    assign data[6128] = ~16'b0;
    assign data[6129] = ~16'b0;
    assign data[6130] = 16'b0;
    assign data[6131] = 16'b0;
    assign data[6132] = ~16'b0;
    assign data[6133] = ~16'b0;
    assign data[6134] = ~16'b0;
    assign data[6135] = ~16'b0;
    assign data[6136] = ~16'b0;
    assign data[6137] = ~16'b0;
    assign data[6138] = ~16'b0;
    assign data[6139] = ~16'b0;
    assign data[6140] = 16'b0;
    assign data[6141] = 16'b0;
    assign data[6142] = ~16'b0;
    assign data[6143] = ~16'b0;
    assign data[6144] = ~16'b0;
    assign data[6145] = ~16'b0;
    assign data[6146] = ~16'b0;
    assign data[6147] = ~16'b0;
    assign data[6148] = ~16'b0;
    assign data[6149] = ~16'b0;
    assign data[6150] = 16'b0;
    assign data[6151] = 16'b0;
    assign data[6152] = ~16'b0;
    assign data[6153] = ~16'b0;
    assign data[6154] = ~16'b0;
    assign data[6155] = ~16'b0;
    assign data[6156] = ~16'b0;
    assign data[6157] = ~16'b0;
    assign data[6158] = ~16'b0;
    assign data[6159] = ~16'b0;
    assign data[6160] = 16'b0;
    assign data[6161] = 16'b0;
    assign data[6162] = 16'b0;
    assign data[6163] = 16'b0;
    assign data[6164] = 16'b0;
    assign data[6165] = 16'b0;
    assign data[6166] = 16'b0;
    assign data[6167] = 16'b0;
    assign data[6168] = 16'b0;
    assign data[6169] = 16'b0;
    assign data[6170] = 16'b0;
    assign data[6171] = 16'b0;
    assign data[6172] = 16'b0;
    assign data[6173] = 16'b0;
    assign data[6174] = 16'b0;
    assign data[6175] = 16'b0;
    assign data[6176] = 16'b0;
    assign data[6177] = 16'b0;
    assign data[6178] = 16'b0;
    assign data[6179] = 16'b0;
    assign data[6180] = ~16'b0;
    assign data[6181] = ~16'b0;
    assign data[6182] = ~16'b0;
    assign data[6183] = ~16'b0;
    assign data[6184] = ~16'b0;
    assign data[6185] = ~16'b0;
    assign data[6186] = ~16'b0;
    assign data[6187] = ~16'b0;
    assign data[6188] = ~16'b0;
    assign data[6189] = ~16'b0;
    assign data[6190] = ~16'b0;
    assign data[6191] = ~16'b0;
    assign data[6192] = ~16'b0;
    assign data[6193] = ~16'b0;
    assign data[6194] = ~16'b0;
    assign data[6195] = ~16'b0;
    assign data[6196] = ~16'b0;
    assign data[6197] = ~16'b0;
    assign data[6198] = ~16'b0;
    assign data[6199] = ~16'b0;
    assign data[6200] = ~16'b0;
    assign data[6201] = ~16'b0;
    assign data[6202] = ~16'b0;
    assign data[6203] = ~16'b0;
    assign data[6204] = ~16'b0;
    assign data[6205] = ~16'b0;
    assign data[6206] = ~16'b0;
    assign data[6207] = ~16'b0;
    assign data[6208] = ~16'b0;
    assign data[6209] = ~16'b0;
    assign data[6210] = ~16'b0;
    assign data[6211] = ~16'b0;
    assign data[6212] = ~16'b0;
    assign data[6213] = ~16'b0;
    assign data[6214] = ~16'b0;
    assign data[6215] = ~16'b0;
    assign data[6216] = ~16'b0;
    assign data[6217] = ~16'b0;
    assign data[6218] = ~16'b0;
    assign data[6219] = ~16'b0;
    assign data[6220] = ~16'b0;
    assign data[6221] = ~16'b0;
    assign data[6222] = ~16'b0;
    assign data[6223] = ~16'b0;
    assign data[6224] = ~16'b0;
    assign data[6225] = ~16'b0;
    assign data[6226] = ~16'b0;
    assign data[6227] = ~16'b0;
    assign data[6228] = ~16'b0;
    assign data[6229] = ~16'b0;
    assign data[6230] = ~16'b0;
    assign data[6231] = ~16'b0;
    assign data[6232] = ~16'b0;
    assign data[6233] = ~16'b0;
    assign data[6234] = ~16'b0;
    assign data[6235] = ~16'b0;
    assign data[6236] = ~16'b0;
    assign data[6237] = ~16'b0;
    assign data[6238] = ~16'b0;
    assign data[6239] = ~16'b0;
    assign data[6240] = ~16'b0;
    assign data[6241] = ~16'b0;
    assign data[6242] = ~16'b0;
    assign data[6243] = ~16'b0;
    assign data[6244] = ~16'b0;
    assign data[6245] = ~16'b0;
    assign data[6246] = ~16'b0;
    assign data[6247] = ~16'b0;
    assign data[6248] = ~16'b0;
    assign data[6249] = ~16'b0;
    assign data[6250] = ~16'b0;
    assign data[6251] = ~16'b0;
    assign data[6252] = ~16'b0;
    assign data[6253] = ~16'b0;
    assign data[6254] = ~16'b0;
    assign data[6255] = ~16'b0;
    assign data[6256] = ~16'b0;
    assign data[6257] = ~16'b0;
    assign data[6258] = ~16'b0;
    assign data[6259] = ~16'b0;
    assign data[6260] = ~16'b0;
    assign data[6261] = ~16'b0;
    assign data[6262] = ~16'b0;
    assign data[6263] = ~16'b0;
    assign data[6264] = ~16'b0;
    assign data[6265] = ~16'b0;
    assign data[6266] = ~16'b0;
    assign data[6267] = ~16'b0;
    assign data[6268] = ~16'b0;
    assign data[6269] = ~16'b0;
    assign data[6270] = ~16'b0;
    assign data[6271] = ~16'b0;
    assign data[6272] = ~16'b0;
    assign data[6273] = ~16'b0;
    assign data[6274] = ~16'b0;
    assign data[6275] = ~16'b0;
    assign data[6276] = ~16'b0;
    assign data[6277] = ~16'b0;
    assign data[6278] = ~16'b0;
    assign data[6279] = ~16'b0;
    assign data[6280] = 16'b0;
    assign data[6281] = 16'b0;
    assign data[6282] = 16'b0;
    assign data[6283] = 16'b0;
    assign data[6284] = 16'b0;
    assign data[6285] = 16'b0;
    assign data[6286] = 16'b0;
    assign data[6287] = 16'b0;
    assign data[6288] = 16'b0;
    assign data[6289] = 16'b0;
    assign data[6290] = 16'b0;
    assign data[6291] = 16'b0;
    assign data[6292] = 16'b0;
    assign data[6293] = 16'b0;
    assign data[6294] = 16'b0;
    assign data[6295] = 16'b0;
    assign data[6296] = 16'b0;
    assign data[6297] = 16'b0;
    assign data[6298] = 16'b0;
    assign data[6299] = 16'b0;
    assign data[6300] = 16'b0;
    assign data[6301] = 16'b0;
    assign data[6302] = ~16'b0;
    assign data[6303] = ~16'b0;
    assign data[6304] = ~16'b0;
    assign data[6305] = ~16'b0;
    assign data[6306] = ~16'b0;
    assign data[6307] = ~16'b0;
    assign data[6308] = ~16'b0;
    assign data[6309] = ~16'b0;
    assign data[6310] = 16'b0;
    assign data[6311] = 16'b0;
    assign data[6312] = ~16'b0;
    assign data[6313] = ~16'b0;
    assign data[6314] = ~16'b0;
    assign data[6315] = ~16'b0;
    assign data[6316] = ~16'b0;
    assign data[6317] = ~16'b0;
    assign data[6318] = ~16'b0;
    assign data[6319] = ~16'b0;
    assign data[6320] = 16'b0;
    assign data[6321] = 16'b0;
    assign data[6322] = ~16'b0;
    assign data[6323] = ~16'b0;
    assign data[6324] = ~16'b0;
    assign data[6325] = ~16'b0;
    assign data[6326] = ~16'b0;
    assign data[6327] = ~16'b0;
    assign data[6328] = ~16'b0;
    assign data[6329] = ~16'b0;
    assign data[6330] = 16'b0;
    assign data[6331] = 16'b0;
    assign data[6332] = ~16'b0;
    assign data[6333] = ~16'b0;
    assign data[6334] = ~16'b0;
    assign data[6335] = ~16'b0;
    assign data[6336] = ~16'b0;
    assign data[6337] = ~16'b0;
    assign data[6338] = ~16'b0;
    assign data[6339] = ~16'b0;
    assign data[6340] = 16'b0;
    assign data[6341] = 16'b0;
    assign data[6342] = ~16'b0;
    assign data[6343] = ~16'b0;
    assign data[6344] = ~16'b0;
    assign data[6345] = ~16'b0;
    assign data[6346] = ~16'b0;
    assign data[6347] = ~16'b0;
    assign data[6348] = ~16'b0;
    assign data[6349] = ~16'b0;
    assign data[6350] = 16'b0;
    assign data[6351] = 16'b0;
    assign data[6352] = ~16'b0;
    assign data[6353] = ~16'b0;
    assign data[6354] = ~16'b0;
    assign data[6355] = ~16'b0;
    assign data[6356] = ~16'b0;
    assign data[6357] = ~16'b0;
    assign data[6358] = ~16'b0;
    assign data[6359] = ~16'b0;
    assign data[6360] = 16'b0;
    assign data[6361] = 16'b0;
    assign data[6362] = ~16'b0;
    assign data[6363] = ~16'b0;
    assign data[6364] = ~16'b0;
    assign data[6365] = ~16'b0;
    assign data[6366] = ~16'b0;
    assign data[6367] = ~16'b0;
    assign data[6368] = ~16'b0;
    assign data[6369] = ~16'b0;
    assign data[6370] = 16'b0;
    assign data[6371] = 16'b0;
    assign data[6372] = ~16'b0;
    assign data[6373] = ~16'b0;
    assign data[6374] = ~16'b0;
    assign data[6375] = ~16'b0;
    assign data[6376] = ~16'b0;
    assign data[6377] = ~16'b0;
    assign data[6378] = ~16'b0;
    assign data[6379] = ~16'b0;
    assign data[6380] = 16'b0;
    assign data[6381] = 16'b0;
    assign data[6382] = ~16'b0;
    assign data[6383] = ~16'b0;
    assign data[6384] = ~16'b0;
    assign data[6385] = ~16'b0;
    assign data[6386] = ~16'b0;
    assign data[6387] = ~16'b0;
    assign data[6388] = ~16'b0;
    assign data[6389] = ~16'b0;
    assign data[6390] = 16'b0;
    assign data[6391] = 16'b0;
    assign data[6392] = ~16'b0;
    assign data[6393] = ~16'b0;
    assign data[6394] = ~16'b0;
    assign data[6395] = ~16'b0;
    assign data[6396] = ~16'b0;
    assign data[6397] = ~16'b0;
    assign data[6398] = ~16'b0;
    assign data[6399] = ~16'b0;
    assign data[6400] = 16'b0;
    assign data[6401] = 16'b0;
    assign data[6402] = ~16'b0;
    assign data[6403] = ~16'b0;
    assign data[6404] = ~16'b0;
    assign data[6405] = ~16'b0;
    assign data[6406] = ~16'b0;
    assign data[6407] = ~16'b0;
    assign data[6408] = ~16'b0;
    assign data[6409] = ~16'b0;
    assign data[6410] = 16'b0;
    assign data[6411] = 16'b0;
    assign data[6412] = ~16'b0;
    assign data[6413] = ~16'b0;
    assign data[6414] = ~16'b0;
    assign data[6415] = ~16'b0;
    assign data[6416] = ~16'b0;
    assign data[6417] = ~16'b0;
    assign data[6418] = ~16'b0;
    assign data[6419] = ~16'b0;
    assign data[6420] = 16'b0;
    assign data[6421] = 16'b0;
    assign data[6422] = ~16'b0;
    assign data[6423] = ~16'b0;
    assign data[6424] = ~16'b0;
    assign data[6425] = ~16'b0;
    assign data[6426] = ~16'b0;
    assign data[6427] = ~16'b0;
    assign data[6428] = ~16'b0;
    assign data[6429] = ~16'b0;
    assign data[6430] = 16'b0;
    assign data[6431] = 16'b0;
    assign data[6432] = ~16'b0;
    assign data[6433] = ~16'b0;
    assign data[6434] = ~16'b0;
    assign data[6435] = ~16'b0;
    assign data[6436] = ~16'b0;
    assign data[6437] = ~16'b0;
    assign data[6438] = ~16'b0;
    assign data[6439] = ~16'b0;
    assign data[6440] = 16'b0;
    assign data[6441] = 16'b0;
    assign data[6442] = ~16'b0;
    assign data[6443] = ~16'b0;
    assign data[6444] = ~16'b0;
    assign data[6445] = ~16'b0;
    assign data[6446] = ~16'b0;
    assign data[6447] = ~16'b0;
    assign data[6448] = ~16'b0;
    assign data[6449] = ~16'b0;
    assign data[6450] = 16'b0;
    assign data[6451] = 16'b0;
    assign data[6452] = ~16'b0;
    assign data[6453] = ~16'b0;
    assign data[6454] = ~16'b0;
    assign data[6455] = ~16'b0;
    assign data[6456] = ~16'b0;
    assign data[6457] = ~16'b0;
    assign data[6458] = ~16'b0;
    assign data[6459] = ~16'b0;
    assign data[6460] = 16'b0;
    assign data[6461] = 16'b0;
    assign data[6462] = ~16'b0;
    assign data[6463] = ~16'b0;
    assign data[6464] = ~16'b0;
    assign data[6465] = ~16'b0;
    assign data[6466] = ~16'b0;
    assign data[6467] = ~16'b0;
    assign data[6468] = ~16'b0;
    assign data[6469] = ~16'b0;
    assign data[6470] = 16'b0;
    assign data[6471] = 16'b0;
    assign data[6472] = ~16'b0;
    assign data[6473] = ~16'b0;
    assign data[6474] = ~16'b0;
    assign data[6475] = ~16'b0;
    assign data[6476] = ~16'b0;
    assign data[6477] = ~16'b0;
    assign data[6478] = ~16'b0;
    assign data[6479] = ~16'b0;
    assign data[6480] = 16'b0;
    assign data[6481] = 16'b0;
    assign data[6482] = ~16'b0;
    assign data[6483] = ~16'b0;
    assign data[6484] = ~16'b0;
    assign data[6485] = ~16'b0;
    assign data[6486] = ~16'b0;
    assign data[6487] = ~16'b0;
    assign data[6488] = ~16'b0;
    assign data[6489] = ~16'b0;
    assign data[6490] = 16'b0;
    assign data[6491] = 16'b0;
    assign data[6492] = ~16'b0;
    assign data[6493] = ~16'b0;
    assign data[6494] = ~16'b0;
    assign data[6495] = ~16'b0;
    assign data[6496] = ~16'b0;
    assign data[6497] = ~16'b0;
    assign data[6498] = ~16'b0;
    assign data[6499] = ~16'b0;
    assign data[6500] = 16'b0;
    assign data[6501] = 16'b0;
    assign data[6502] = ~16'b0;
    assign data[6503] = ~16'b0;
    assign data[6504] = ~16'b0;
    assign data[6505] = ~16'b0;
    assign data[6506] = ~16'b0;
    assign data[6507] = ~16'b0;
    assign data[6508] = ~16'b0;
    assign data[6509] = ~16'b0;
    assign data[6510] = 16'b0;
    assign data[6511] = 16'b0;
    assign data[6512] = ~16'b0;
    assign data[6513] = ~16'b0;
    assign data[6514] = ~16'b0;
    assign data[6515] = ~16'b0;
    assign data[6516] = ~16'b0;
    assign data[6517] = ~16'b0;
    assign data[6518] = ~16'b0;
    assign data[6519] = ~16'b0;
    assign data[6520] = 16'b0;
    assign data[6521] = 16'b0;
    assign data[6522] = ~16'b0;
    assign data[6523] = ~16'b0;
    assign data[6524] = ~16'b0;
    assign data[6525] = ~16'b0;
    assign data[6526] = ~16'b0;
    assign data[6527] = ~16'b0;
    assign data[6528] = ~16'b0;
    assign data[6529] = ~16'b0;
    assign data[6530] = 16'b0;
    assign data[6531] = 16'b0;
    assign data[6532] = ~16'b0;
    assign data[6533] = ~16'b0;
    assign data[6534] = ~16'b0;
    assign data[6535] = ~16'b0;
    assign data[6536] = ~16'b0;
    assign data[6537] = ~16'b0;
    assign data[6538] = ~16'b0;
    assign data[6539] = ~16'b0;
    assign data[6540] = 16'b0;
    assign data[6541] = 16'b0;
    assign data[6542] = ~16'b0;
    assign data[6543] = ~16'b0;
    assign data[6544] = ~16'b0;
    assign data[6545] = ~16'b0;
    assign data[6546] = ~16'b0;
    assign data[6547] = ~16'b0;
    assign data[6548] = ~16'b0;
    assign data[6549] = ~16'b0;
    assign data[6550] = 16'b0;
    assign data[6551] = 16'b0;
    assign data[6552] = ~16'b0;
    assign data[6553] = ~16'b0;
    assign data[6554] = ~16'b0;
    assign data[6555] = ~16'b0;
    assign data[6556] = ~16'b0;
    assign data[6557] = ~16'b0;
    assign data[6558] = ~16'b0;
    assign data[6559] = ~16'b0;
    assign data[6560] = 16'b0;
    assign data[6561] = 16'b0;
    assign data[6562] = ~16'b0;
    assign data[6563] = ~16'b0;
    assign data[6564] = ~16'b0;
    assign data[6565] = ~16'b0;
    assign data[6566] = ~16'b0;
    assign data[6567] = ~16'b0;
    assign data[6568] = ~16'b0;
    assign data[6569] = ~16'b0;
    assign data[6570] = 16'b0;
    assign data[6571] = 16'b0;
    assign data[6572] = ~16'b0;
    assign data[6573] = ~16'b0;
    assign data[6574] = ~16'b0;
    assign data[6575] = ~16'b0;
    assign data[6576] = ~16'b0;
    assign data[6577] = ~16'b0;
    assign data[6578] = ~16'b0;
    assign data[6579] = ~16'b0;
    assign data[6580] = 16'b0;
    assign data[6581] = 16'b0;
    assign data[6582] = ~16'b0;
    assign data[6583] = ~16'b0;
    assign data[6584] = ~16'b0;
    assign data[6585] = ~16'b0;
    assign data[6586] = ~16'b0;
    assign data[6587] = ~16'b0;
    assign data[6588] = ~16'b0;
    assign data[6589] = ~16'b0;
    assign data[6590] = 16'b0;
    assign data[6591] = 16'b0;
    assign data[6592] = ~16'b0;
    assign data[6593] = ~16'b0;
    assign data[6594] = ~16'b0;
    assign data[6595] = ~16'b0;
    assign data[6596] = ~16'b0;
    assign data[6597] = ~16'b0;
    assign data[6598] = ~16'b0;
    assign data[6599] = ~16'b0;
    assign data[6600] = 16'b0;
    assign data[6601] = 16'b0;
    assign data[6602] = ~16'b0;
    assign data[6603] = ~16'b0;
    assign data[6604] = ~16'b0;
    assign data[6605] = ~16'b0;
    assign data[6606] = ~16'b0;
    assign data[6607] = ~16'b0;
    assign data[6608] = ~16'b0;
    assign data[6609] = ~16'b0;
    assign data[6610] = 16'b0;
    assign data[6611] = 16'b0;
    assign data[6612] = ~16'b0;
    assign data[6613] = ~16'b0;
    assign data[6614] = ~16'b0;
    assign data[6615] = ~16'b0;
    assign data[6616] = ~16'b0;
    assign data[6617] = ~16'b0;
    assign data[6618] = ~16'b0;
    assign data[6619] = ~16'b0;
    assign data[6620] = 16'b0;
    assign data[6621] = 16'b0;
    assign data[6622] = ~16'b0;
    assign data[6623] = ~16'b0;
    assign data[6624] = ~16'b0;
    assign data[6625] = ~16'b0;
    assign data[6626] = ~16'b0;
    assign data[6627] = ~16'b0;
    assign data[6628] = ~16'b0;
    assign data[6629] = ~16'b0;
    assign data[6630] = 16'b0;
    assign data[6631] = 16'b0;
    assign data[6632] = ~16'b0;
    assign data[6633] = ~16'b0;
    assign data[6634] = ~16'b0;
    assign data[6635] = ~16'b0;
    assign data[6636] = ~16'b0;
    assign data[6637] = ~16'b0;
    assign data[6638] = ~16'b0;
    assign data[6639] = ~16'b0;
    assign data[6640] = 16'b0;
    assign data[6641] = 16'b0;
    assign data[6642] = ~16'b0;
    assign data[6643] = ~16'b0;
    assign data[6644] = ~16'b0;
    assign data[6645] = ~16'b0;
    assign data[6646] = ~16'b0;
    assign data[6647] = ~16'b0;
    assign data[6648] = ~16'b0;
    assign data[6649] = ~16'b0;
    assign data[6650] = 16'b0;
    assign data[6651] = 16'b0;
    assign data[6652] = ~16'b0;
    assign data[6653] = ~16'b0;
    assign data[6654] = ~16'b0;
    assign data[6655] = ~16'b0;
    assign data[6656] = ~16'b0;
    assign data[6657] = ~16'b0;
    assign data[6658] = ~16'b0;
    assign data[6659] = ~16'b0;
    assign data[6660] = 16'b0;
    assign data[6661] = 16'b0;
    assign data[6662] = 16'b0;
    assign data[6663] = 16'b0;
    assign data[6664] = 16'b0;
    assign data[6665] = 16'b0;
    assign data[6666] = 16'b0;
    assign data[6667] = 16'b0;
    assign data[6668] = 16'b0;
    assign data[6669] = 16'b0;
    assign data[6670] = 16'b0;
    assign data[6671] = 16'b0;
    assign data[6672] = 16'b0;
    assign data[6673] = 16'b0;
    assign data[6674] = 16'b0;
    assign data[6675] = 16'b0;
    assign data[6676] = 16'b0;
    assign data[6677] = 16'b0;
    assign data[6678] = 16'b0;
    assign data[6679] = 16'b0;
    assign data[6680] = ~16'b0;
    assign data[6681] = ~16'b0;
    assign data[6682] = ~16'b0;
    assign data[6683] = ~16'b0;
    assign data[6684] = ~16'b0;
    assign data[6685] = ~16'b0;
    assign data[6686] = ~16'b0;
    assign data[6687] = ~16'b0;
    assign data[6688] = ~16'b0;
    assign data[6689] = ~16'b0;
    assign data[6690] = ~16'b0;
    assign data[6691] = ~16'b0;
    assign data[6692] = ~16'b0;
    assign data[6693] = ~16'b0;
    assign data[6694] = ~16'b0;
    assign data[6695] = ~16'b0;
    assign data[6696] = ~16'b0;
    assign data[6697] = ~16'b0;
    assign data[6698] = ~16'b0;
    assign data[6699] = ~16'b0;
    assign data[6700] = ~16'b0;
    assign data[6701] = ~16'b0;
    assign data[6702] = ~16'b0;
    assign data[6703] = ~16'b0;
    assign data[6704] = ~16'b0;
    assign data[6705] = ~16'b0;
    assign data[6706] = ~16'b0;
    assign data[6707] = ~16'b0;
    assign data[6708] = ~16'b0;
    assign data[6709] = ~16'b0;
    assign data[6710] = ~16'b0;
    assign data[6711] = ~16'b0;
    assign data[6712] = ~16'b0;
    assign data[6713] = ~16'b0;
    assign data[6714] = ~16'b0;
    assign data[6715] = ~16'b0;
    assign data[6716] = ~16'b0;
    assign data[6717] = ~16'b0;
    assign data[6718] = ~16'b0;
    assign data[6719] = ~16'b0;
    assign data[6720] = ~16'b0;
    assign data[6721] = ~16'b0;
    assign data[6722] = ~16'b0;
    assign data[6723] = ~16'b0;
    assign data[6724] = ~16'b0;
    assign data[6725] = ~16'b0;
    assign data[6726] = ~16'b0;
    assign data[6727] = ~16'b0;
    assign data[6728] = ~16'b0;
    assign data[6729] = ~16'b0;
    assign data[6730] = ~16'b0;
    assign data[6731] = ~16'b0;
    assign data[6732] = ~16'b0;
    assign data[6733] = ~16'b0;
    assign data[6734] = ~16'b0;
    assign data[6735] = ~16'b0;
    assign data[6736] = ~16'b0;
    assign data[6737] = ~16'b0;
    assign data[6738] = ~16'b0;
    assign data[6739] = ~16'b0;
    assign data[6740] = ~16'b0;
    assign data[6741] = ~16'b0;
    assign data[6742] = ~16'b0;
    assign data[6743] = ~16'b0;
    assign data[6744] = ~16'b0;
    assign data[6745] = ~16'b0;
    assign data[6746] = ~16'b0;
    assign data[6747] = ~16'b0;
    assign data[6748] = ~16'b0;
    assign data[6749] = ~16'b0;
    assign data[6750] = ~16'b0;
    assign data[6751] = ~16'b0;
    assign data[6752] = ~16'b0;
    assign data[6753] = ~16'b0;
    assign data[6754] = ~16'b0;
    assign data[6755] = ~16'b0;
    assign data[6756] = ~16'b0;
    assign data[6757] = ~16'b0;
    assign data[6758] = ~16'b0;
    assign data[6759] = ~16'b0;
    assign data[6760] = ~16'b0;
    assign data[6761] = ~16'b0;
    assign data[6762] = ~16'b0;
    assign data[6763] = ~16'b0;
    assign data[6764] = ~16'b0;
    assign data[6765] = ~16'b0;
    assign data[6766] = ~16'b0;
    assign data[6767] = ~16'b0;
    assign data[6768] = ~16'b0;
    assign data[6769] = ~16'b0;
    assign data[6770] = ~16'b0;
    assign data[6771] = ~16'b0;
    assign data[6772] = ~16'b0;
    assign data[6773] = ~16'b0;
    assign data[6774] = ~16'b0;
    assign data[6775] = ~16'b0;
    assign data[6776] = ~16'b0;
    assign data[6777] = ~16'b0;
    assign data[6778] = ~16'b0;
    assign data[6779] = ~16'b0;
    assign data[6780] = ~16'b0;
    assign data[6781] = ~16'b0;
    assign data[6782] = ~16'b0;
    assign data[6783] = ~16'b0;
    assign data[6784] = ~16'b0;
    assign data[6785] = ~16'b0;
    assign data[6786] = ~16'b0;
    assign data[6787] = ~16'b0;
    assign data[6788] = ~16'b0;
    assign data[6789] = ~16'b0;
    assign data[6790] = ~16'b0;
    assign data[6791] = ~16'b0;
    assign data[6792] = ~16'b0;
    assign data[6793] = ~16'b0;
    assign data[6794] = ~16'b0;
    assign data[6795] = ~16'b0;
    assign data[6796] = ~16'b0;
    assign data[6797] = ~16'b0;
    assign data[6798] = ~16'b0;
    assign data[6799] = ~16'b0;
    assign data[6800] = ~16'b0;
    assign data[6801] = ~16'b0;
    assign data[6802] = ~16'b0;
    assign data[6803] = ~16'b0;
    assign data[6804] = ~16'b0;
    assign data[6805] = ~16'b0;
    assign data[6806] = ~16'b0;
    assign data[6807] = ~16'b0;
    assign data[6808] = ~16'b0;
    assign data[6809] = ~16'b0;
    assign data[6810] = ~16'b0;
    assign data[6811] = ~16'b0;
    assign data[6812] = ~16'b0;
    assign data[6813] = ~16'b0;
    assign data[6814] = ~16'b0;
    assign data[6815] = ~16'b0;
    assign data[6816] = ~16'b0;
    assign data[6817] = ~16'b0;
    assign data[6818] = ~16'b0;
    assign data[6819] = ~16'b0;
    assign data[6820] = ~16'b0;
    assign data[6821] = ~16'b0;
    assign data[6822] = ~16'b0;
    assign data[6823] = ~16'b0;
    assign data[6824] = ~16'b0;
    assign data[6825] = ~16'b0;
    assign data[6826] = ~16'b0;
    assign data[6827] = ~16'b0;
    assign data[6828] = ~16'b0;
    assign data[6829] = ~16'b0;
    assign data[6830] = ~16'b0;
    assign data[6831] = ~16'b0;
    assign data[6832] = ~16'b0;
    assign data[6833] = ~16'b0;
    assign data[6834] = ~16'b0;
    assign data[6835] = ~16'b0;
    assign data[6836] = ~16'b0;
    assign data[6837] = ~16'b0;
    assign data[6838] = ~16'b0;
    assign data[6839] = ~16'b0;
    assign data[6840] = ~16'b0;
    assign data[6841] = ~16'b0;
    assign data[6842] = ~16'b0;
    assign data[6843] = ~16'b0;
    assign data[6844] = ~16'b0;
    assign data[6845] = ~16'b0;
    assign data[6846] = ~16'b0;
    assign data[6847] = ~16'b0;
    assign data[6848] = ~16'b0;
    assign data[6849] = ~16'b0;
    assign data[6850] = 16'b0;
    assign data[6851] = 16'b0;
    assign data[6852] = 16'b0;
    assign data[6853] = 16'b0;
    assign data[6854] = 16'b0;
    assign data[6855] = 16'b0;
    assign data[6856] = 16'b0;
    assign data[6857] = 16'b0;
    assign data[6858] = 16'b0;
    assign data[6859] = 16'b0;
    assign data[6860] = 16'b0;
    assign data[6861] = 16'b0;
    assign data[6862] = 16'b0;
    assign data[6863] = 16'b0;
    assign data[6864] = 16'b0;
    assign data[6865] = 16'b0;
    assign data[6866] = 16'b0;
    assign data[6867] = 16'b0;
    assign data[6868] = 16'b0;
    assign data[6869] = 16'b0;
    assign data[6870] = 16'b0;
    assign data[6871] = 16'b0;
    assign data[6872] = ~16'b0;
    assign data[6873] = ~16'b0;
    assign data[6874] = ~16'b0;
    assign data[6875] = ~16'b0;
    assign data[6876] = ~16'b0;
    assign data[6877] = ~16'b0;
    assign data[6878] = ~16'b0;
    assign data[6879] = ~16'b0;
    assign data[6880] = 16'b0;
    assign data[6881] = 16'b0;
    assign data[6882] = ~16'b0;
    assign data[6883] = ~16'b0;
    assign data[6884] = ~16'b0;
    assign data[6885] = ~16'b0;
    assign data[6886] = ~16'b0;
    assign data[6887] = ~16'b0;
    assign data[6888] = ~16'b0;
    assign data[6889] = ~16'b0;
    assign data[6890] = 16'b0;
    assign data[6891] = 16'b0;
    assign data[6892] = ~16'b0;
    assign data[6893] = ~16'b0;
    assign data[6894] = ~16'b0;
    assign data[6895] = ~16'b0;
    assign data[6896] = ~16'b0;
    assign data[6897] = ~16'b0;
    assign data[6898] = ~16'b0;
    assign data[6899] = ~16'b0;
    assign data[6900] = 16'b0;
    assign data[6901] = 16'b0;
    assign data[6902] = ~16'b0;
    assign data[6903] = ~16'b0;
    assign data[6904] = ~16'b0;
    assign data[6905] = ~16'b0;
    assign data[6906] = ~16'b0;
    assign data[6907] = ~16'b0;
    assign data[6908] = ~16'b0;
    assign data[6909] = ~16'b0;
    assign data[6910] = 16'b0;
    assign data[6911] = 16'b0;
    assign data[6912] = ~16'b0;
    assign data[6913] = ~16'b0;
    assign data[6914] = ~16'b0;
    assign data[6915] = ~16'b0;
    assign data[6916] = ~16'b0;
    assign data[6917] = ~16'b0;
    assign data[6918] = ~16'b0;
    assign data[6919] = ~16'b0;
    assign data[6920] = 16'b0;
    assign data[6921] = 16'b0;
    assign data[6922] = ~16'b0;
    assign data[6923] = ~16'b0;
    assign data[6924] = ~16'b0;
    assign data[6925] = ~16'b0;
    assign data[6926] = ~16'b0;
    assign data[6927] = ~16'b0;
    assign data[6928] = ~16'b0;
    assign data[6929] = ~16'b0;
    assign data[6930] = 16'b0;
    assign data[6931] = 16'b0;
    assign data[6932] = ~16'b0;
    assign data[6933] = ~16'b0;
    assign data[6934] = ~16'b0;
    assign data[6935] = ~16'b0;
    assign data[6936] = ~16'b0;
    assign data[6937] = ~16'b0;
    assign data[6938] = ~16'b0;
    assign data[6939] = ~16'b0;
    assign data[6940] = 16'b0;
    assign data[6941] = 16'b0;
    assign data[6942] = ~16'b0;
    assign data[6943] = ~16'b0;
    assign data[6944] = ~16'b0;
    assign data[6945] = ~16'b0;
    assign data[6946] = ~16'b0;
    assign data[6947] = ~16'b0;
    assign data[6948] = ~16'b0;
    assign data[6949] = ~16'b0;
    assign data[6950] = 16'b0;
    assign data[6951] = 16'b0;
    assign data[6952] = ~16'b0;
    assign data[6953] = ~16'b0;
    assign data[6954] = ~16'b0;
    assign data[6955] = ~16'b0;
    assign data[6956] = ~16'b0;
    assign data[6957] = ~16'b0;
    assign data[6958] = ~16'b0;
    assign data[6959] = ~16'b0;
    assign data[6960] = 16'b0;
    assign data[6961] = 16'b0;
    assign data[6962] = ~16'b0;
    assign data[6963] = ~16'b0;
    assign data[6964] = ~16'b0;
    assign data[6965] = ~16'b0;
    assign data[6966] = ~16'b0;
    assign data[6967] = ~16'b0;
    assign data[6968] = ~16'b0;
    assign data[6969] = ~16'b0;
    assign data[6970] = 16'b0;
    assign data[6971] = 16'b0;
    assign data[6972] = ~16'b0;
    assign data[6973] = ~16'b0;
    assign data[6974] = ~16'b0;
    assign data[6975] = ~16'b0;
    assign data[6976] = ~16'b0;
    assign data[6977] = ~16'b0;
    assign data[6978] = ~16'b0;
    assign data[6979] = ~16'b0;
    assign data[6980] = 16'b0;
    assign data[6981] = 16'b0;
    assign data[6982] = ~16'b0;
    assign data[6983] = ~16'b0;
    assign data[6984] = ~16'b0;
    assign data[6985] = ~16'b0;
    assign data[6986] = ~16'b0;
    assign data[6987] = ~16'b0;
    assign data[6988] = ~16'b0;
    assign data[6989] = ~16'b0;
    assign data[6990] = 16'b0;
    assign data[6991] = 16'b0;
    assign data[6992] = ~16'b0;
    assign data[6993] = ~16'b0;
    assign data[6994] = ~16'b0;
    assign data[6995] = ~16'b0;
    assign data[6996] = ~16'b0;
    assign data[6997] = ~16'b0;
    assign data[6998] = ~16'b0;
    assign data[6999] = ~16'b0;
    assign data[7000] = 16'b0;
    assign data[7001] = 16'b0;
    assign data[7002] = ~16'b0;
    assign data[7003] = ~16'b0;
    assign data[7004] = ~16'b0;
    assign data[7005] = ~16'b0;
    assign data[7006] = ~16'b0;
    assign data[7007] = ~16'b0;
    assign data[7008] = ~16'b0;
    assign data[7009] = ~16'b0;
    assign data[7010] = 16'b0;
    assign data[7011] = 16'b0;
    assign data[7012] = ~16'b0;
    assign data[7013] = ~16'b0;
    assign data[7014] = ~16'b0;
    assign data[7015] = ~16'b0;
    assign data[7016] = ~16'b0;
    assign data[7017] = ~16'b0;
    assign data[7018] = ~16'b0;
    assign data[7019] = ~16'b0;
    assign data[7020] = 16'b0;
    assign data[7021] = 16'b0;
    assign data[7022] = ~16'b0;
    assign data[7023] = ~16'b0;
    assign data[7024] = ~16'b0;
    assign data[7025] = ~16'b0;
    assign data[7026] = ~16'b0;
    assign data[7027] = ~16'b0;
    assign data[7028] = ~16'b0;
    assign data[7029] = ~16'b0;
    assign data[7030] = 16'b0;
    assign data[7031] = 16'b0;
    assign data[7032] = ~16'b0;
    assign data[7033] = ~16'b0;
    assign data[7034] = ~16'b0;
    assign data[7035] = ~16'b0;
    assign data[7036] = ~16'b0;
    assign data[7037] = ~16'b0;
    assign data[7038] = ~16'b0;
    assign data[7039] = ~16'b0;
    assign data[7040] = 16'b0;
    assign data[7041] = 16'b0;
    assign data[7042] = ~16'b0;
    assign data[7043] = ~16'b0;
    assign data[7044] = ~16'b0;
    assign data[7045] = ~16'b0;
    assign data[7046] = ~16'b0;
    assign data[7047] = ~16'b0;
    assign data[7048] = ~16'b0;
    assign data[7049] = ~16'b0;
    assign data[7050] = 16'b0;
    assign data[7051] = 16'b0;
    assign data[7052] = ~16'b0;
    assign data[7053] = ~16'b0;
    assign data[7054] = ~16'b0;
    assign data[7055] = ~16'b0;
    assign data[7056] = ~16'b0;
    assign data[7057] = ~16'b0;
    assign data[7058] = ~16'b0;
    assign data[7059] = ~16'b0;
    assign data[7060] = 16'b0;
    assign data[7061] = 16'b0;
    assign data[7062] = ~16'b0;
    assign data[7063] = ~16'b0;
    assign data[7064] = ~16'b0;
    assign data[7065] = ~16'b0;
    assign data[7066] = ~16'b0;
    assign data[7067] = ~16'b0;
    assign data[7068] = ~16'b0;
    assign data[7069] = ~16'b0;
    assign data[7070] = 16'b0;
    assign data[7071] = 16'b0;
    assign data[7072] = ~16'b0;
    assign data[7073] = ~16'b0;
    assign data[7074] = ~16'b0;
    assign data[7075] = ~16'b0;
    assign data[7076] = ~16'b0;
    assign data[7077] = ~16'b0;
    assign data[7078] = ~16'b0;
    assign data[7079] = ~16'b0;
    assign data[7080] = 16'b0;
    assign data[7081] = 16'b0;
    assign data[7082] = 16'b0;
    assign data[7083] = 16'b0;
    assign data[7084] = 16'b0;
    assign data[7085] = 16'b0;
    assign data[7086] = 16'b0;
    assign data[7087] = 16'b0;
    assign data[7088] = 16'b0;
    assign data[7089] = 16'b0;
    assign data[7090] = 16'b0;
    assign data[7091] = 16'b0;
    assign data[7092] = 16'b0;
    assign data[7093] = 16'b0;
    assign data[7094] = 16'b0;
    assign data[7095] = 16'b0;
    assign data[7096] = 16'b0;
    assign data[7097] = 16'b0;
    assign data[7098] = 16'b0;
    assign data[7099] = 16'b0;
    assign data[7100] = ~16'b0;
    assign data[7101] = ~16'b0;
    assign data[7102] = ~16'b0;
    assign data[7103] = ~16'b0;
    assign data[7104] = ~16'b0;
    assign data[7105] = ~16'b0;
    assign data[7106] = ~16'b0;
    assign data[7107] = ~16'b0;
    assign data[7108] = ~16'b0;
    assign data[7109] = ~16'b0;
    assign data[7110] = ~16'b0;
    assign data[7111] = ~16'b0;
    assign data[7112] = ~16'b0;
    assign data[7113] = ~16'b0;
    assign data[7114] = ~16'b0;
    assign data[7115] = ~16'b0;
    assign data[7116] = ~16'b0;
    assign data[7117] = ~16'b0;
    assign data[7118] = ~16'b0;
    assign data[7119] = ~16'b0;
    assign data[7120] = ~16'b0;
    assign data[7121] = ~16'b0;
    assign data[7122] = ~16'b0;
    assign data[7123] = ~16'b0;
    assign data[7124] = ~16'b0;
    assign data[7125] = ~16'b0;
    assign data[7126] = ~16'b0;
    assign data[7127] = ~16'b0;
    assign data[7128] = ~16'b0;
    assign data[7129] = ~16'b0;
    assign data[7130] = ~16'b0;
    assign data[7131] = ~16'b0;
    assign data[7132] = ~16'b0;
    assign data[7133] = ~16'b0;
    assign data[7134] = ~16'b0;
    assign data[7135] = ~16'b0;
    assign data[7136] = ~16'b0;
    assign data[7137] = ~16'b0;
    assign data[7138] = ~16'b0;
    assign data[7139] = ~16'b0;
    assign data[7140] = ~16'b0;
    assign data[7141] = ~16'b0;
    assign data[7142] = ~16'b0;
    assign data[7143] = ~16'b0;
    assign data[7144] = ~16'b0;
    assign data[7145] = ~16'b0;
    assign data[7146] = ~16'b0;
    assign data[7147] = ~16'b0;
    assign data[7148] = ~16'b0;
    assign data[7149] = ~16'b0;
    assign data[7150] = ~16'b0;
    assign data[7151] = ~16'b0;
    assign data[7152] = ~16'b0;
    assign data[7153] = ~16'b0;
    assign data[7154] = ~16'b0;
    assign data[7155] = ~16'b0;
    assign data[7156] = ~16'b0;
    assign data[7157] = ~16'b0;
    assign data[7158] = ~16'b0;
    assign data[7159] = ~16'b0;
    assign data[7160] = ~16'b0;
    assign data[7161] = ~16'b0;
    assign data[7162] = ~16'b0;
    assign data[7163] = ~16'b0;
    assign data[7164] = ~16'b0;
    assign data[7165] = ~16'b0;
    assign data[7166] = ~16'b0;
    assign data[7167] = ~16'b0;
    assign data[7168] = ~16'b0;
    assign data[7169] = ~16'b0;
    assign data[7170] = ~16'b0;
    assign data[7171] = ~16'b0;
    assign data[7172] = ~16'b0;
    assign data[7173] = ~16'b0;
    assign data[7174] = ~16'b0;
    assign data[7175] = ~16'b0;
    assign data[7176] = ~16'b0;
    assign data[7177] = ~16'b0;
    assign data[7178] = ~16'b0;
    assign data[7179] = ~16'b0;
    assign data[7180] = ~16'b0;
    assign data[7181] = ~16'b0;
    assign data[7182] = ~16'b0;
    assign data[7183] = ~16'b0;
    assign data[7184] = ~16'b0;
    assign data[7185] = ~16'b0;
    assign data[7186] = ~16'b0;
    assign data[7187] = ~16'b0;
    assign data[7188] = ~16'b0;
    assign data[7189] = ~16'b0;
    assign data[7190] = ~16'b0;
    assign data[7191] = ~16'b0;
    assign data[7192] = ~16'b0;
    assign data[7193] = ~16'b0;
    assign data[7194] = ~16'b0;
    assign data[7195] = ~16'b0;
    assign data[7196] = ~16'b0;
    assign data[7197] = ~16'b0;
    assign data[7198] = ~16'b0;
    assign data[7199] = ~16'b0;
    assign data[7200] = ~16'b0;
    assign data[7201] = ~16'b0;
    assign data[7202] = ~16'b0;
    assign data[7203] = ~16'b0;
    assign data[7204] = ~16'b0;
    assign data[7205] = ~16'b0;
    assign data[7206] = ~16'b0;
    assign data[7207] = ~16'b0;
    assign data[7208] = ~16'b0;
    assign data[7209] = ~16'b0;
    assign data[7210] = ~16'b0;
    assign data[7211] = ~16'b0;
    assign data[7212] = ~16'b0;
    assign data[7213] = ~16'b0;
    assign data[7214] = ~16'b0;
    assign data[7215] = ~16'b0;
    assign data[7216] = ~16'b0;
    assign data[7217] = ~16'b0;
    assign data[7218] = ~16'b0;
    assign data[7219] = ~16'b0;
    assign data[7220] = 16'b0;
    assign data[7221] = 16'b0;
    assign data[7222] = 16'b0;
    assign data[7223] = 16'b0;
    assign data[7224] = 16'b0;
    assign data[7225] = 16'b0;
    assign data[7226] = 16'b0;
    assign data[7227] = 16'b0;
    assign data[7228] = 16'b0;
    assign data[7229] = 16'b0;
    assign data[7230] = 16'b0;
    assign data[7231] = 16'b0;
    assign data[7232] = 16'b0;
    assign data[7233] = 16'b0;
    assign data[7234] = 16'b0;
    assign data[7235] = 16'b0;
    assign data[7236] = 16'b0;
    assign data[7237] = 16'b0;
    assign data[7238] = 16'b0;
    assign data[7239] = 16'b0;
    assign data[7240] = 16'b0;
    assign data[7241] = 16'b0;
    assign data[7242] = ~16'b0;
    assign data[7243] = ~16'b0;
    assign data[7244] = ~16'b0;
    assign data[7245] = ~16'b0;
    assign data[7246] = ~16'b0;
    assign data[7247] = ~16'b0;
    assign data[7248] = ~16'b0;
    assign data[7249] = ~16'b0;
    assign data[7250] = 16'b0;
    assign data[7251] = 16'b0;
    assign data[7252] = ~16'b0;
    assign data[7253] = ~16'b0;
    assign data[7254] = ~16'b0;
    assign data[7255] = ~16'b0;
    assign data[7256] = ~16'b0;
    assign data[7257] = ~16'b0;
    assign data[7258] = ~16'b0;
    assign data[7259] = ~16'b0;
    assign data[7260] = 16'b0;
    assign data[7261] = 16'b0;
    assign data[7262] = ~16'b0;
    assign data[7263] = ~16'b0;
    assign data[7264] = ~16'b0;
    assign data[7265] = ~16'b0;
    assign data[7266] = ~16'b0;
    assign data[7267] = ~16'b0;
    assign data[7268] = ~16'b0;
    assign data[7269] = ~16'b0;
    assign data[7270] = 16'b0;
    assign data[7271] = 16'b0;
    assign data[7272] = ~16'b0;
    assign data[7273] = ~16'b0;
    assign data[7274] = ~16'b0;
    assign data[7275] = ~16'b0;
    assign data[7276] = ~16'b0;
    assign data[7277] = ~16'b0;
    assign data[7278] = ~16'b0;
    assign data[7279] = ~16'b0;
    assign data[7280] = 16'b0;
    assign data[7281] = 16'b0;
    assign data[7282] = ~16'b0;
    assign data[7283] = ~16'b0;
    assign data[7284] = ~16'b0;
    assign data[7285] = ~16'b0;
    assign data[7286] = ~16'b0;
    assign data[7287] = ~16'b0;
    assign data[7288] = ~16'b0;
    assign data[7289] = ~16'b0;
    assign data[7290] = 16'b0;
    assign data[7291] = 16'b0;
    assign data[7292] = ~16'b0;
    assign data[7293] = ~16'b0;
    assign data[7294] = ~16'b0;
    assign data[7295] = ~16'b0;
    assign data[7296] = ~16'b0;
    assign data[7297] = ~16'b0;
    assign data[7298] = ~16'b0;
    assign data[7299] = ~16'b0;
    assign data[7300] = 16'b0;
    assign data[7301] = 16'b0;
    assign data[7302] = ~16'b0;
    assign data[7303] = ~16'b0;
    assign data[7304] = ~16'b0;
    assign data[7305] = ~16'b0;
    assign data[7306] = ~16'b0;
    assign data[7307] = ~16'b0;
    assign data[7308] = ~16'b0;
    assign data[7309] = ~16'b0;
    assign data[7310] = 16'b0;
    assign data[7311] = 16'b0;
    assign data[7312] = ~16'b0;
    assign data[7313] = ~16'b0;
    assign data[7314] = ~16'b0;
    assign data[7315] = ~16'b0;
    assign data[7316] = ~16'b0;
    assign data[7317] = ~16'b0;
    assign data[7318] = ~16'b0;
    assign data[7319] = ~16'b0;
    assign data[7320] = 16'b0;
    assign data[7321] = 16'b0;
    assign data[7322] = ~16'b0;
    assign data[7323] = ~16'b0;
    assign data[7324] = ~16'b0;
    assign data[7325] = ~16'b0;
    assign data[7326] = ~16'b0;
    assign data[7327] = ~16'b0;
    assign data[7328] = ~16'b0;
    assign data[7329] = ~16'b0;
    assign data[7330] = 16'b0;
    assign data[7331] = 16'b0;
    assign data[7332] = ~16'b0;
    assign data[7333] = ~16'b0;
    assign data[7334] = ~16'b0;
    assign data[7335] = ~16'b0;
    assign data[7336] = ~16'b0;
    assign data[7337] = ~16'b0;
    assign data[7338] = ~16'b0;
    assign data[7339] = ~16'b0;
    assign data[7340] = 16'b0;
    assign data[7341] = 16'b0;
    assign data[7342] = ~16'b0;
    assign data[7343] = ~16'b0;
    assign data[7344] = ~16'b0;
    assign data[7345] = ~16'b0;
    assign data[7346] = ~16'b0;
    assign data[7347] = ~16'b0;
    assign data[7348] = ~16'b0;
    assign data[7349] = ~16'b0;
    assign data[7350] = 16'b0;
    assign data[7351] = 16'b0;
    assign data[7352] = ~16'b0;
    assign data[7353] = ~16'b0;
    assign data[7354] = ~16'b0;
    assign data[7355] = ~16'b0;
    assign data[7356] = ~16'b0;
    assign data[7357] = ~16'b0;
    assign data[7358] = ~16'b0;
    assign data[7359] = ~16'b0;
    assign data[7360] = 16'b0;
    assign data[7361] = 16'b0;
    assign data[7362] = ~16'b0;
    assign data[7363] = ~16'b0;
    assign data[7364] = ~16'b0;
    assign data[7365] = ~16'b0;
    assign data[7366] = ~16'b0;
    assign data[7367] = ~16'b0;
    assign data[7368] = ~16'b0;
    assign data[7369] = ~16'b0;
    assign data[7370] = 16'b0;
    assign data[7371] = 16'b0;
    assign data[7372] = ~16'b0;
    assign data[7373] = ~16'b0;
    assign data[7374] = ~16'b0;
    assign data[7375] = ~16'b0;
    assign data[7376] = ~16'b0;
    assign data[7377] = ~16'b0;
    assign data[7378] = ~16'b0;
    assign data[7379] = ~16'b0;
    assign data[7380] = 16'b0;
    assign data[7381] = 16'b0;
    assign data[7382] = ~16'b0;
    assign data[7383] = ~16'b0;
    assign data[7384] = ~16'b0;
    assign data[7385] = ~16'b0;
    assign data[7386] = ~16'b0;
    assign data[7387] = ~16'b0;
    assign data[7388] = ~16'b0;
    assign data[7389] = ~16'b0;
    assign data[7390] = 16'b0;
    assign data[7391] = 16'b0;
    assign data[7392] = ~16'b0;
    assign data[7393] = ~16'b0;
    assign data[7394] = ~16'b0;
    assign data[7395] = ~16'b0;
    assign data[7396] = ~16'b0;
    assign data[7397] = ~16'b0;
    assign data[7398] = ~16'b0;
    assign data[7399] = ~16'b0;
    assign data[7400] = 16'b0;
    assign data[7401] = 16'b0;
    assign data[7402] = 16'b0;
    assign data[7403] = 16'b0;
    assign data[7404] = 16'b0;
    assign data[7405] = 16'b0;
    assign data[7406] = 16'b0;
    assign data[7407] = 16'b0;
    assign data[7408] = 16'b0;
    assign data[7409] = 16'b0;
    assign data[7410] = 16'b0;
    assign data[7411] = 16'b0;
    assign data[7412] = 16'b0;
    assign data[7413] = 16'b0;
    assign data[7414] = 16'b0;
    assign data[7415] = 16'b0;
    assign data[7416] = 16'b0;
    assign data[7417] = 16'b0;
    assign data[7418] = 16'b0;
    assign data[7419] = 16'b0;
    assign data[7420] = ~16'b0;
    assign data[7421] = ~16'b0;
    assign data[7422] = ~16'b0;
    assign data[7423] = ~16'b0;
    assign data[7424] = ~16'b0;
    assign data[7425] = ~16'b0;
    assign data[7426] = ~16'b0;
    assign data[7427] = ~16'b0;
    assign data[7428] = ~16'b0;
    assign data[7429] = ~16'b0;
    assign data[7430] = ~16'b0;
    assign data[7431] = ~16'b0;
    assign data[7432] = ~16'b0;
    assign data[7433] = ~16'b0;
    assign data[7434] = ~16'b0;
    assign data[7435] = ~16'b0;
    assign data[7436] = ~16'b0;
    assign data[7437] = ~16'b0;
    assign data[7438] = ~16'b0;
    assign data[7439] = ~16'b0;
    assign data[7440] = ~16'b0;
    assign data[7441] = ~16'b0;
    assign data[7442] = ~16'b0;
    assign data[7443] = ~16'b0;
    assign data[7444] = ~16'b0;
    assign data[7445] = ~16'b0;
    assign data[7446] = ~16'b0;
    assign data[7447] = ~16'b0;
    assign data[7448] = ~16'b0;
    assign data[7449] = ~16'b0;
    assign data[7450] = ~16'b0;
    assign data[7451] = ~16'b0;
    assign data[7452] = ~16'b0;
    assign data[7453] = ~16'b0;
    assign data[7454] = ~16'b0;
    assign data[7455] = ~16'b0;
    assign data[7456] = ~16'b0;
    assign data[7457] = ~16'b0;
    assign data[7458] = ~16'b0;
    assign data[7459] = ~16'b0;
    assign data[7460] = ~16'b0;
    assign data[7461] = ~16'b0;
    assign data[7462] = ~16'b0;
    assign data[7463] = ~16'b0;
    assign data[7464] = ~16'b0;
    assign data[7465] = ~16'b0;
    assign data[7466] = ~16'b0;
    assign data[7467] = ~16'b0;
    assign data[7468] = ~16'b0;
    assign data[7469] = ~16'b0;
    assign data[7470] = ~16'b0;
    assign data[7471] = ~16'b0;
    assign data[7472] = ~16'b0;
    assign data[7473] = ~16'b0;
    assign data[7474] = ~16'b0;
    assign data[7475] = ~16'b0;
    assign data[7476] = ~16'b0;
    assign data[7477] = ~16'b0;
    assign data[7478] = ~16'b0;
    assign data[7479] = ~16'b0;
    assign data[7480] = ~16'b0;
    assign data[7481] = ~16'b0;
    assign data[7482] = ~16'b0;
    assign data[7483] = ~16'b0;
    assign data[7484] = ~16'b0;
    assign data[7485] = ~16'b0;
    assign data[7486] = ~16'b0;
    assign data[7487] = ~16'b0;
    assign data[7488] = ~16'b0;
    assign data[7489] = ~16'b0;
    assign data[7490] = ~16'b0;
    assign data[7491] = ~16'b0;
    assign data[7492] = ~16'b0;
    assign data[7493] = ~16'b0;
    assign data[7494] = ~16'b0;
    assign data[7495] = ~16'b0;
    assign data[7496] = ~16'b0;
    assign data[7497] = ~16'b0;
    assign data[7498] = ~16'b0;
    assign data[7499] = ~16'b0;
    assign data[7500] = ~16'b0;
    assign data[7501] = ~16'b0;
    assign data[7502] = ~16'b0;
    assign data[7503] = ~16'b0;
    assign data[7504] = ~16'b0;
    assign data[7505] = ~16'b0;
    assign data[7506] = ~16'b0;
    assign data[7507] = ~16'b0;
    assign data[7508] = ~16'b0;
    assign data[7509] = ~16'b0;
    assign data[7510] = ~16'b0;
    assign data[7511] = ~16'b0;
    assign data[7512] = ~16'b0;
    assign data[7513] = ~16'b0;
    assign data[7514] = ~16'b0;
    assign data[7515] = ~16'b0;
    assign data[7516] = ~16'b0;
    assign data[7517] = ~16'b0;
    assign data[7518] = ~16'b0;
    assign data[7519] = ~16'b0;
    assign data[7520] = ~16'b0;
    assign data[7521] = ~16'b0;
    assign data[7522] = ~16'b0;
    assign data[7523] = ~16'b0;
    assign data[7524] = ~16'b0;
    assign data[7525] = ~16'b0;
    assign data[7526] = ~16'b0;
    assign data[7527] = ~16'b0;
    assign data[7528] = ~16'b0;
    assign data[7529] = ~16'b0;
    assign data[7530] = ~16'b0;
    assign data[7531] = ~16'b0;
    assign data[7532] = ~16'b0;
    assign data[7533] = ~16'b0;
    assign data[7534] = ~16'b0;
    assign data[7535] = ~16'b0;
    assign data[7536] = ~16'b0;
    assign data[7537] = ~16'b0;
    assign data[7538] = ~16'b0;
    assign data[7539] = ~16'b0;
    assign data[7540] = ~16'b0;
    assign data[7541] = ~16'b0;
    assign data[7542] = ~16'b0;
    assign data[7543] = ~16'b0;
    assign data[7544] = ~16'b0;
    assign data[7545] = ~16'b0;
    assign data[7546] = ~16'b0;
    assign data[7547] = ~16'b0;
    assign data[7548] = ~16'b0;
    assign data[7549] = ~16'b0;
    assign data[7550] = 16'b0;
    assign data[7551] = 16'b0;
    assign data[7552] = 16'b0;
    assign data[7553] = 16'b0;
    assign data[7554] = 16'b0;
    assign data[7555] = 16'b0;
    assign data[7556] = 16'b0;
    assign data[7557] = 16'b0;
    assign data[7558] = 16'b0;
    assign data[7559] = 16'b0;
    assign data[7560] = 16'b0;
    assign data[7561] = 16'b0;
    assign data[7562] = 16'b0;
    assign data[7563] = 16'b0;
    assign data[7564] = 16'b0;
    assign data[7565] = 16'b0;
    assign data[7566] = 16'b0;
    assign data[7567] = 16'b0;
    assign data[7568] = 16'b0;
    assign data[7569] = 16'b0;
    assign data[7570] = 16'b0;
    assign data[7571] = 16'b0;
    assign data[7572] = ~16'b0;
    assign data[7573] = ~16'b0;
    assign data[7574] = ~16'b0;
    assign data[7575] = ~16'b0;
    assign data[7576] = ~16'b0;
    assign data[7577] = ~16'b0;
    assign data[7578] = ~16'b0;
    assign data[7579] = ~16'b0;
    assign data[7580] = 16'b0;
    assign data[7581] = 16'b0;
    assign data[7582] = ~16'b0;
    assign data[7583] = ~16'b0;
    assign data[7584] = ~16'b0;
    assign data[7585] = ~16'b0;
    assign data[7586] = ~16'b0;
    assign data[7587] = ~16'b0;
    assign data[7588] = ~16'b0;
    assign data[7589] = ~16'b0;
    assign data[7590] = 16'b0;
    assign data[7591] = 16'b0;
    assign data[7592] = ~16'b0;
    assign data[7593] = ~16'b0;
    assign data[7594] = ~16'b0;
    assign data[7595] = ~16'b0;
    assign data[7596] = ~16'b0;
    assign data[7597] = ~16'b0;
    assign data[7598] = ~16'b0;
    assign data[7599] = ~16'b0;
    assign data[7600] = 16'b0;
    assign data[7601] = 16'b0;
    assign data[7602] = ~16'b0;
    assign data[7603] = ~16'b0;
    assign data[7604] = ~16'b0;
    assign data[7605] = ~16'b0;
    assign data[7606] = ~16'b0;
    assign data[7607] = ~16'b0;
    assign data[7608] = ~16'b0;
    assign data[7609] = ~16'b0;
    assign data[7610] = 16'b0;
    assign data[7611] = 16'b0;
    assign data[7612] = ~16'b0;
    assign data[7613] = ~16'b0;
    assign data[7614] = ~16'b0;
    assign data[7615] = ~16'b0;
    assign data[7616] = ~16'b0;
    assign data[7617] = ~16'b0;
    assign data[7618] = ~16'b0;
    assign data[7619] = ~16'b0;
    assign data[7620] = 16'b0;
    assign data[7621] = 16'b0;
    assign data[7622] = ~16'b0;
    assign data[7623] = ~16'b0;
    assign data[7624] = ~16'b0;
    assign data[7625] = ~16'b0;
    assign data[7626] = ~16'b0;
    assign data[7627] = ~16'b0;
    assign data[7628] = ~16'b0;
    assign data[7629] = ~16'b0;
    assign data[7630] = 16'b0;
    assign data[7631] = 16'b0;
    assign data[7632] = ~16'b0;
    assign data[7633] = ~16'b0;
    assign data[7634] = ~16'b0;
    assign data[7635] = ~16'b0;
    assign data[7636] = ~16'b0;
    assign data[7637] = ~16'b0;
    assign data[7638] = ~16'b0;
    assign data[7639] = ~16'b0;
    assign data[7640] = 16'b0;
    assign data[7641] = 16'b0;
    assign data[7642] = ~16'b0;
    assign data[7643] = ~16'b0;
    assign data[7644] = ~16'b0;
    assign data[7645] = ~16'b0;
    assign data[7646] = ~16'b0;
    assign data[7647] = ~16'b0;
    assign data[7648] = ~16'b0;
    assign data[7649] = ~16'b0;
    assign data[7650] = 16'b0;
    assign data[7651] = 16'b0;
    assign data[7652] = ~16'b0;
    assign data[7653] = ~16'b0;
    assign data[7654] = ~16'b0;
    assign data[7655] = ~16'b0;
    assign data[7656] = ~16'b0;
    assign data[7657] = ~16'b0;
    assign data[7658] = ~16'b0;
    assign data[7659] = ~16'b0;
    assign data[7660] = 16'b0;
    assign data[7661] = 16'b0;
    assign data[7662] = ~16'b0;
    assign data[7663] = ~16'b0;
    assign data[7664] = ~16'b0;
    assign data[7665] = ~16'b0;
    assign data[7666] = ~16'b0;
    assign data[7667] = ~16'b0;
    assign data[7668] = ~16'b0;
    assign data[7669] = ~16'b0;
    assign data[7670] = 16'b0;
    assign data[7671] = 16'b0;
    assign data[7672] = ~16'b0;
    assign data[7673] = ~16'b0;
    assign data[7674] = ~16'b0;
    assign data[7675] = ~16'b0;
    assign data[7676] = ~16'b0;
    assign data[7677] = ~16'b0;
    assign data[7678] = ~16'b0;
    assign data[7679] = ~16'b0;
    assign data[7680] = 16'b0;
    assign data[7681] = 16'b0;
    assign data[7682] = ~16'b0;
    assign data[7683] = ~16'b0;
    assign data[7684] = ~16'b0;
    assign data[7685] = ~16'b0;
    assign data[7686] = ~16'b0;
    assign data[7687] = ~16'b0;
    assign data[7688] = ~16'b0;
    assign data[7689] = ~16'b0;
    assign data[7690] = 16'b0;
    assign data[7691] = 16'b0;
    assign data[7692] = ~16'b0;
    assign data[7693] = ~16'b0;
    assign data[7694] = ~16'b0;
    assign data[7695] = ~16'b0;
    assign data[7696] = ~16'b0;
    assign data[7697] = ~16'b0;
    assign data[7698] = ~16'b0;
    assign data[7699] = ~16'b0;
    assign data[7700] = 16'b0;
    assign data[7701] = 16'b0;
    assign data[7702] = ~16'b0;
    assign data[7703] = ~16'b0;
    assign data[7704] = ~16'b0;
    assign data[7705] = ~16'b0;
    assign data[7706] = ~16'b0;
    assign data[7707] = ~16'b0;
    assign data[7708] = ~16'b0;
    assign data[7709] = ~16'b0;
    assign data[7710] = 16'b0;
    assign data[7711] = 16'b0;
    assign data[7712] = ~16'b0;
    assign data[7713] = ~16'b0;
    assign data[7714] = ~16'b0;
    assign data[7715] = ~16'b0;
    assign data[7716] = ~16'b0;
    assign data[7717] = ~16'b0;
    assign data[7718] = ~16'b0;
    assign data[7719] = ~16'b0;
    assign data[7720] = 16'b0;
    assign data[7721] = 16'b0;
    assign data[7722] = ~16'b0;
    assign data[7723] = ~16'b0;
    assign data[7724] = ~16'b0;
    assign data[7725] = ~16'b0;
    assign data[7726] = ~16'b0;
    assign data[7727] = ~16'b0;
    assign data[7728] = ~16'b0;
    assign data[7729] = ~16'b0;
    assign data[7730] = 16'b0;
    assign data[7731] = 16'b0;
    assign data[7732] = ~16'b0;
    assign data[7733] = ~16'b0;
    assign data[7734] = ~16'b0;
    assign data[7735] = ~16'b0;
    assign data[7736] = ~16'b0;
    assign data[7737] = ~16'b0;
    assign data[7738] = ~16'b0;
    assign data[7739] = ~16'b0;
    assign data[7740] = 16'b0;
    assign data[7741] = 16'b0;
    assign data[7742] = ~16'b0;
    assign data[7743] = ~16'b0;
    assign data[7744] = ~16'b0;
    assign data[7745] = ~16'b0;
    assign data[7746] = ~16'b0;
    assign data[7747] = ~16'b0;
    assign data[7748] = ~16'b0;
    assign data[7749] = ~16'b0;
    assign data[7750] = 16'b0;
    assign data[7751] = 16'b0;
    assign data[7752] = ~16'b0;
    assign data[7753] = ~16'b0;
    assign data[7754] = ~16'b0;
    assign data[7755] = ~16'b0;
    assign data[7756] = ~16'b0;
    assign data[7757] = ~16'b0;
    assign data[7758] = ~16'b0;
    assign data[7759] = ~16'b0;
    assign data[7760] = 16'b0;
    assign data[7761] = 16'b0;
    assign data[7762] = ~16'b0;
    assign data[7763] = ~16'b0;
    assign data[7764] = ~16'b0;
    assign data[7765] = ~16'b0;
    assign data[7766] = ~16'b0;
    assign data[7767] = ~16'b0;
    assign data[7768] = ~16'b0;
    assign data[7769] = ~16'b0;
    assign data[7770] = 16'b0;
    assign data[7771] = 16'b0;
    assign data[7772] = ~16'b0;
    assign data[7773] = ~16'b0;
    assign data[7774] = ~16'b0;
    assign data[7775] = ~16'b0;
    assign data[7776] = ~16'b0;
    assign data[7777] = ~16'b0;
    assign data[7778] = ~16'b0;
    assign data[7779] = ~16'b0;
    assign data[7780] = 16'b0;
    assign data[7781] = 16'b0;
    assign data[7782] = ~16'b0;
    assign data[7783] = ~16'b0;
    assign data[7784] = ~16'b0;
    assign data[7785] = ~16'b0;
    assign data[7786] = ~16'b0;
    assign data[7787] = ~16'b0;
    assign data[7788] = ~16'b0;
    assign data[7789] = ~16'b0;
    assign data[7790] = 16'b0;
    assign data[7791] = 16'b0;
    assign data[7792] = ~16'b0;
    assign data[7793] = ~16'b0;
    assign data[7794] = ~16'b0;
    assign data[7795] = ~16'b0;
    assign data[7796] = ~16'b0;
    assign data[7797] = ~16'b0;
    assign data[7798] = ~16'b0;
    assign data[7799] = ~16'b0;
    assign data[7800] = 16'b0;
    assign data[7801] = 16'b0;
    assign data[7802] = ~16'b0;
    assign data[7803] = ~16'b0;
    assign data[7804] = ~16'b0;
    assign data[7805] = ~16'b0;
    assign data[7806] = ~16'b0;
    assign data[7807] = ~16'b0;
    assign data[7808] = ~16'b0;
    assign data[7809] = ~16'b0;
    assign data[7810] = 16'b0;
    assign data[7811] = 16'b0;
    assign data[7812] = ~16'b0;
    assign data[7813] = ~16'b0;
    assign data[7814] = ~16'b0;
    assign data[7815] = ~16'b0;
    assign data[7816] = ~16'b0;
    assign data[7817] = ~16'b0;
    assign data[7818] = ~16'b0;
    assign data[7819] = ~16'b0;
    assign data[7820] = 16'b0;
    assign data[7821] = 16'b0;
    assign data[7822] = ~16'b0;
    assign data[7823] = ~16'b0;
    assign data[7824] = ~16'b0;
    assign data[7825] = ~16'b0;
    assign data[7826] = ~16'b0;
    assign data[7827] = ~16'b0;
    assign data[7828] = ~16'b0;
    assign data[7829] = ~16'b0;
    assign data[7830] = 16'b0;
    assign data[7831] = 16'b0;
    assign data[7832] = ~16'b0;
    assign data[7833] = ~16'b0;
    assign data[7834] = ~16'b0;
    assign data[7835] = ~16'b0;
    assign data[7836] = ~16'b0;
    assign data[7837] = ~16'b0;
    assign data[7838] = ~16'b0;
    assign data[7839] = ~16'b0;
    assign data[7840] = 16'b0;
    assign data[7841] = 16'b0;
    assign data[7842] = ~16'b0;
    assign data[7843] = ~16'b0;
    assign data[7844] = ~16'b0;
    assign data[7845] = ~16'b0;
    assign data[7846] = ~16'b0;
    assign data[7847] = ~16'b0;
    assign data[7848] = ~16'b0;
    assign data[7849] = ~16'b0;
    assign data[7850] = 16'b0;
    assign data[7851] = 16'b0;
    assign data[7852] = ~16'b0;
    assign data[7853] = ~16'b0;
    assign data[7854] = ~16'b0;
    assign data[7855] = ~16'b0;
    assign data[7856] = ~16'b0;
    assign data[7857] = ~16'b0;
    assign data[7858] = ~16'b0;
    assign data[7859] = ~16'b0;
    assign data[7860] = 16'b0;
    assign data[7861] = 16'b0;
    assign data[7862] = 16'b0;
    assign data[7863] = 16'b0;
    assign data[7864] = 16'b0;
    assign data[7865] = 16'b0;
    assign data[7866] = 16'b0;
    assign data[7867] = 16'b0;
    assign data[7868] = 16'b0;
    assign data[7869] = 16'b0;
    assign data[7870] = 16'b0;
    assign data[7871] = 16'b0;
    assign data[7872] = 16'b0;
    assign data[7873] = 16'b0;
    assign data[7874] = 16'b0;
    assign data[7875] = 16'b0;
    assign data[7876] = 16'b0;
    assign data[7877] = 16'b0;
    assign data[7878] = 16'b0;
    assign data[7879] = 16'b0;
    assign data[7880] = ~16'b0;
    assign data[7881] = ~16'b0;
    assign data[7882] = ~16'b0;
    assign data[7883] = ~16'b0;
    assign data[7884] = ~16'b0;
    assign data[7885] = ~16'b0;
    assign data[7886] = ~16'b0;
    assign data[7887] = ~16'b0;
    assign data[7888] = ~16'b0;
    assign data[7889] = ~16'b0;
    assign data[7890] = ~16'b0;
    assign data[7891] = ~16'b0;
    assign data[7892] = ~16'b0;
    assign data[7893] = ~16'b0;
    assign data[7894] = ~16'b0;
    assign data[7895] = ~16'b0;
    assign data[7896] = ~16'b0;
    assign data[7897] = ~16'b0;
    assign data[7898] = ~16'b0;
    assign data[7899] = ~16'b0;
    assign data[7900] = ~16'b0;
    assign data[7901] = ~16'b0;
    assign data[7902] = ~16'b0;
    assign data[7903] = ~16'b0;
    assign data[7904] = ~16'b0;
    assign data[7905] = ~16'b0;
    assign data[7906] = ~16'b0;
    assign data[7907] = ~16'b0;
    assign data[7908] = ~16'b0;
    assign data[7909] = ~16'b0;
    assign data[7910] = ~16'b0;
    assign data[7911] = ~16'b0;
    assign data[7912] = ~16'b0;
    assign data[7913] = ~16'b0;
    assign data[7914] = ~16'b0;
    assign data[7915] = ~16'b0;
    assign data[7916] = ~16'b0;
    assign data[7917] = ~16'b0;
    assign data[7918] = ~16'b0;
    assign data[7919] = ~16'b0;
    assign data[7920] = ~16'b0;
    assign data[7921] = ~16'b0;
    assign data[7922] = ~16'b0;
    assign data[7923] = ~16'b0;
    assign data[7924] = ~16'b0;
    assign data[7925] = ~16'b0;
    assign data[7926] = ~16'b0;
    assign data[7927] = ~16'b0;
    assign data[7928] = ~16'b0;
    assign data[7929] = ~16'b0;
    assign data[7930] = ~16'b0;
    assign data[7931] = ~16'b0;
    assign data[7932] = ~16'b0;
    assign data[7933] = ~16'b0;
    assign data[7934] = ~16'b0;
    assign data[7935] = ~16'b0;
    assign data[7936] = ~16'b0;
    assign data[7937] = ~16'b0;
    assign data[7938] = ~16'b0;
    assign data[7939] = ~16'b0;
    assign data[7940] = ~16'b0;
    assign data[7941] = ~16'b0;
    assign data[7942] = ~16'b0;
    assign data[7943] = ~16'b0;
    assign data[7944] = ~16'b0;
    assign data[7945] = ~16'b0;
    assign data[7946] = ~16'b0;
    assign data[7947] = ~16'b0;
    assign data[7948] = ~16'b0;
    assign data[7949] = ~16'b0;
    assign data[7950] = ~16'b0;
    assign data[7951] = ~16'b0;
    assign data[7952] = ~16'b0;
    assign data[7953] = ~16'b0;
    assign data[7954] = ~16'b0;
    assign data[7955] = ~16'b0;
    assign data[7956] = ~16'b0;
    assign data[7957] = ~16'b0;
    assign data[7958] = ~16'b0;
    assign data[7959] = ~16'b0;
    assign data[7960] = ~16'b0;
    assign data[7961] = ~16'b0;
    assign data[7962] = ~16'b0;
    assign data[7963] = ~16'b0;
    assign data[7964] = ~16'b0;
    assign data[7965] = ~16'b0;
    assign data[7966] = ~16'b0;
    assign data[7967] = ~16'b0;
    assign data[7968] = ~16'b0;
    assign data[7969] = ~16'b0;
    assign data[7970] = ~16'b0;
    assign data[7971] = ~16'b0;
    assign data[7972] = ~16'b0;
    assign data[7973] = ~16'b0;
    assign data[7974] = ~16'b0;
    assign data[7975] = ~16'b0;
    assign data[7976] = ~16'b0;
    assign data[7977] = ~16'b0;
    assign data[7978] = ~16'b0;
    assign data[7979] = ~16'b0;
    assign data[7980] = ~16'b0;
    assign data[7981] = ~16'b0;
    assign data[7982] = ~16'b0;
    assign data[7983] = ~16'b0;
    assign data[7984] = ~16'b0;
    assign data[7985] = ~16'b0;
    assign data[7986] = ~16'b0;
    assign data[7987] = ~16'b0;
    assign data[7988] = ~16'b0;
    assign data[7989] = ~16'b0;
    assign data[7990] = ~16'b0;
    assign data[7991] = ~16'b0;
    assign data[7992] = ~16'b0;
    assign data[7993] = ~16'b0;
    assign data[7994] = ~16'b0;
    assign data[7995] = ~16'b0;
    assign data[7996] = ~16'b0;
    assign data[7997] = ~16'b0;
    assign data[7998] = ~16'b0;
    assign data[7999] = ~16'b0;
    assign data[8000] = ~16'b0;
    assign data[8001] = ~16'b0;
    assign data[8002] = ~16'b0;
    assign data[8003] = ~16'b0;
    assign data[8004] = ~16'b0;
    assign data[8005] = ~16'b0;
    assign data[8006] = ~16'b0;
    assign data[8007] = ~16'b0;
    assign data[8008] = ~16'b0;
    assign data[8009] = ~16'b0;
    assign data[8010] = ~16'b0;
    assign data[8011] = ~16'b0;
    assign data[8012] = ~16'b0;
    assign data[8013] = ~16'b0;
    assign data[8014] = ~16'b0;
    assign data[8015] = ~16'b0;
    assign data[8016] = ~16'b0;
    assign data[8017] = ~16'b0;
    assign data[8018] = ~16'b0;
    assign data[8019] = ~16'b0;
    assign data[8020] = ~16'b0;
    assign data[8021] = ~16'b0;
    assign data[8022] = ~16'b0;
    assign data[8023] = ~16'b0;
    assign data[8024] = ~16'b0;
    assign data[8025] = ~16'b0;
    assign data[8026] = ~16'b0;
    assign data[8027] = ~16'b0;
    assign data[8028] = ~16'b0;
    assign data[8029] = ~16'b0;
    assign data[8030] = ~16'b0;
    assign data[8031] = ~16'b0;
    assign data[8032] = ~16'b0;
    assign data[8033] = ~16'b0;
    assign data[8034] = ~16'b0;
    assign data[8035] = ~16'b0;
    assign data[8036] = ~16'b0;
    assign data[8037] = ~16'b0;
    assign data[8038] = ~16'b0;
    assign data[8039] = ~16'b0;
    assign data[8040] = ~16'b0;
    assign data[8041] = ~16'b0;
    assign data[8042] = ~16'b0;
    assign data[8043] = ~16'b0;
    assign data[8044] = ~16'b0;
    assign data[8045] = ~16'b0;
    assign data[8046] = ~16'b0;
    assign data[8047] = ~16'b0;
    assign data[8048] = ~16'b0;
    assign data[8049] = ~16'b0;
    assign data[8050] = ~16'b0;
    assign data[8051] = ~16'b0;
    assign data[8052] = ~16'b0;
    assign data[8053] = ~16'b0;
    assign data[8054] = ~16'b0;
    assign data[8055] = ~16'b0;
    assign data[8056] = ~16'b0;
    assign data[8057] = ~16'b0;
    assign data[8058] = ~16'b0;
    assign data[8059] = ~16'b0;
    assign data[8060] = ~16'b0;
    assign data[8061] = ~16'b0;
    assign data[8062] = ~16'b0;
    assign data[8063] = ~16'b0;
    assign data[8064] = ~16'b0;
    assign data[8065] = ~16'b0;
    assign data[8066] = ~16'b0;
    assign data[8067] = ~16'b0;
    assign data[8068] = ~16'b0;
    assign data[8069] = ~16'b0;
    assign data[8070] = ~16'b0;
    assign data[8071] = ~16'b0;
    assign data[8072] = ~16'b0;
    assign data[8073] = ~16'b0;
    assign data[8074] = ~16'b0;
    assign data[8075] = ~16'b0;
    assign data[8076] = ~16'b0;
    assign data[8077] = ~16'b0;
    assign data[8078] = ~16'b0;
    assign data[8079] = ~16'b0;
    assign data[8080] = ~16'b0;
    assign data[8081] = ~16'b0;
    assign data[8082] = ~16'b0;
    assign data[8083] = ~16'b0;
    assign data[8084] = ~16'b0;
    assign data[8085] = ~16'b0;
    assign data[8086] = ~16'b0;
    assign data[8087] = ~16'b0;
    assign data[8088] = ~16'b0;
    assign data[8089] = ~16'b0;
    assign data[8090] = ~16'b0;
    assign data[8091] = ~16'b0;
    assign data[8092] = ~16'b0;
    assign data[8093] = ~16'b0;
    assign data[8094] = ~16'b0;
    assign data[8095] = ~16'b0;
    assign data[8096] = ~16'b0;
    assign data[8097] = ~16'b0;
    assign data[8098] = ~16'b0;
    assign data[8099] = ~16'b0;
    assign data[8100] = ~16'b0;
    assign data[8101] = ~16'b0;
    assign data[8102] = ~16'b0;
    assign data[8103] = ~16'b0;
    assign data[8104] = ~16'b0;
    assign data[8105] = ~16'b0;
    assign data[8106] = ~16'b0;
    assign data[8107] = ~16'b0;
    assign data[8108] = ~16'b0;
    assign data[8109] = ~16'b0;
    assign data[8110] = ~16'b0;
    assign data[8111] = ~16'b0;
    assign data[8112] = ~16'b0;
    assign data[8113] = ~16'b0;
    assign data[8114] = ~16'b0;
    assign data[8115] = ~16'b0;
    assign data[8116] = ~16'b0;
    assign data[8117] = ~16'b0;
    assign data[8118] = ~16'b0;
    assign data[8119] = ~16'b0;
    assign data[8120] = ~16'b0;
    assign data[8121] = ~16'b0;
    assign data[8122] = ~16'b0;
    assign data[8123] = ~16'b0;
    assign data[8124] = ~16'b0;
    assign data[8125] = ~16'b0;
    assign data[8126] = ~16'b0;
    assign data[8127] = ~16'b0;
    assign data[8128] = ~16'b0;
    assign data[8129] = ~16'b0;
    assign data[8130] = 16'b0;
    assign data[8131] = 16'b0;
    assign data[8132] = 16'b0;
    assign data[8133] = 16'b0;
    assign data[8134] = 16'b0;
    assign data[8135] = 16'b0;
    assign data[8136] = 16'b0;
    assign data[8137] = 16'b0;
    assign data[8138] = 16'b0;
    assign data[8139] = 16'b0;
    assign data[8140] = 16'b0;
    assign data[8141] = 16'b0;
    assign data[8142] = 16'b0;
    assign data[8143] = 16'b0;
    assign data[8144] = 16'b0;
    assign data[8145] = 16'b0;
    assign data[8146] = 16'b0;
    assign data[8147] = 16'b0;
    assign data[8148] = 16'b0;
    assign data[8149] = 16'b0;
    assign data[8150] = 16'b0;
    assign data[8151] = 16'b0;
    assign data[8152] = ~16'b0;
    assign data[8153] = ~16'b0;
    assign data[8154] = ~16'b0;
    assign data[8155] = ~16'b0;
    assign data[8156] = ~16'b0;
    assign data[8157] = ~16'b0;
    assign data[8158] = ~16'b0;
    assign data[8159] = ~16'b0;
    assign data[8160] = 16'b0;
    assign data[8161] = 16'b0;
    assign data[8162] = ~16'b0;
    assign data[8163] = ~16'b0;
    assign data[8164] = ~16'b0;
    assign data[8165] = ~16'b0;
    assign data[8166] = ~16'b0;
    assign data[8167] = ~16'b0;
    assign data[8168] = ~16'b0;
    assign data[8169] = ~16'b0;
    assign data[8170] = 16'b0;
    assign data[8171] = 16'b0;
    assign data[8172] = ~16'b0;
    assign data[8173] = ~16'b0;
    assign data[8174] = ~16'b0;
    assign data[8175] = ~16'b0;
    assign data[8176] = ~16'b0;
    assign data[8177] = ~16'b0;
    assign data[8178] = ~16'b0;
    assign data[8179] = ~16'b0;
    assign data[8180] = 16'b0;
    assign data[8181] = 16'b0;
    assign data[8182] = ~16'b0;
    assign data[8183] = ~16'b0;
    assign data[8184] = ~16'b0;
    assign data[8185] = ~16'b0;
    assign data[8186] = ~16'b0;
    assign data[8187] = ~16'b0;
    assign data[8188] = ~16'b0;
    assign data[8189] = ~16'b0;
    assign data[8190] = 16'b0;
    assign data[8191] = 16'b0;
    assign data[8192] = ~16'b0;
    assign data[8193] = ~16'b0;
    assign data[8194] = ~16'b0;
    assign data[8195] = ~16'b0;
    assign data[8196] = ~16'b0;
    assign data[8197] = ~16'b0;
    assign data[8198] = ~16'b0;
    assign data[8199] = ~16'b0;
    assign data[8200] = 16'b0;
    assign data[8201] = 16'b0;
    assign data[8202] = ~16'b0;
    assign data[8203] = ~16'b0;
    assign data[8204] = ~16'b0;
    assign data[8205] = ~16'b0;
    assign data[8206] = ~16'b0;
    assign data[8207] = ~16'b0;
    assign data[8208] = ~16'b0;
    assign data[8209] = ~16'b0;
    assign data[8210] = 16'b0;
    assign data[8211] = 16'b0;
    assign data[8212] = ~16'b0;
    assign data[8213] = ~16'b0;
    assign data[8214] = ~16'b0;
    assign data[8215] = ~16'b0;
    assign data[8216] = ~16'b0;
    assign data[8217] = ~16'b0;
    assign data[8218] = ~16'b0;
    assign data[8219] = ~16'b0;
    assign data[8220] = 16'b0;
    assign data[8221] = 16'b0;
    assign data[8222] = ~16'b0;
    assign data[8223] = ~16'b0;
    assign data[8224] = ~16'b0;
    assign data[8225] = ~16'b0;
    assign data[8226] = ~16'b0;
    assign data[8227] = ~16'b0;
    assign data[8228] = ~16'b0;
    assign data[8229] = ~16'b0;
    assign data[8230] = 16'b0;
    assign data[8231] = 16'b0;
    assign data[8232] = ~16'b0;
    assign data[8233] = ~16'b0;
    assign data[8234] = ~16'b0;
    assign data[8235] = ~16'b0;
    assign data[8236] = ~16'b0;
    assign data[8237] = ~16'b0;
    assign data[8238] = ~16'b0;
    assign data[8239] = ~16'b0;
    assign data[8240] = 16'b0;
    assign data[8241] = 16'b0;
    assign data[8242] = ~16'b0;
    assign data[8243] = ~16'b0;
    assign data[8244] = ~16'b0;
    assign data[8245] = ~16'b0;
    assign data[8246] = ~16'b0;
    assign data[8247] = ~16'b0;
    assign data[8248] = ~16'b0;
    assign data[8249] = ~16'b0;
    assign data[8250] = 16'b0;
    assign data[8251] = 16'b0;
    assign data[8252] = ~16'b0;
    assign data[8253] = ~16'b0;
    assign data[8254] = ~16'b0;
    assign data[8255] = ~16'b0;
    assign data[8256] = ~16'b0;
    assign data[8257] = ~16'b0;
    assign data[8258] = ~16'b0;
    assign data[8259] = ~16'b0;
    assign data[8260] = 16'b0;
    assign data[8261] = 16'b0;
    assign data[8262] = ~16'b0;
    assign data[8263] = ~16'b0;
    assign data[8264] = ~16'b0;
    assign data[8265] = ~16'b0;
    assign data[8266] = ~16'b0;
    assign data[8267] = ~16'b0;
    assign data[8268] = ~16'b0;
    assign data[8269] = ~16'b0;
    assign data[8270] = 16'b0;
    assign data[8271] = 16'b0;
    assign data[8272] = ~16'b0;
    assign data[8273] = ~16'b0;
    assign data[8274] = ~16'b0;
    assign data[8275] = ~16'b0;
    assign data[8276] = ~16'b0;
    assign data[8277] = ~16'b0;
    assign data[8278] = ~16'b0;
    assign data[8279] = ~16'b0;
    assign data[8280] = 16'b0;
    assign data[8281] = 16'b0;
    assign data[8282] = ~16'b0;
    assign data[8283] = ~16'b0;
    assign data[8284] = ~16'b0;
    assign data[8285] = ~16'b0;
    assign data[8286] = ~16'b0;
    assign data[8287] = ~16'b0;
    assign data[8288] = ~16'b0;
    assign data[8289] = ~16'b0;
    assign data[8290] = 16'b0;
    assign data[8291] = 16'b0;
    assign data[8292] = ~16'b0;
    assign data[8293] = ~16'b0;
    assign data[8294] = ~16'b0;
    assign data[8295] = ~16'b0;
    assign data[8296] = ~16'b0;
    assign data[8297] = ~16'b0;
    assign data[8298] = ~16'b0;
    assign data[8299] = ~16'b0;
    assign data[8300] = 16'b0;
    assign data[8301] = 16'b0;
    assign data[8302] = ~16'b0;
    assign data[8303] = ~16'b0;
    assign data[8304] = ~16'b0;
    assign data[8305] = ~16'b0;
    assign data[8306] = ~16'b0;
    assign data[8307] = ~16'b0;
    assign data[8308] = ~16'b0;
    assign data[8309] = ~16'b0;
    assign data[8310] = 16'b0;
    assign data[8311] = 16'b0;
    assign data[8312] = 16'b0;
    assign data[8313] = 16'b0;
    assign data[8314] = 16'b0;
    assign data[8315] = 16'b0;
    assign data[8316] = 16'b0;
    assign data[8317] = 16'b0;
    assign data[8318] = 16'b0;
    assign data[8319] = 16'b0;
    assign data[8320] = 16'b0;
    assign data[8321] = 16'b0;
    assign data[8322] = 16'b0;
    assign data[8323] = 16'b0;
    assign data[8324] = 16'b0;
    assign data[8325] = 16'b0;
    assign data[8326] = 16'b0;
    assign data[8327] = 16'b0;
    assign data[8328] = 16'b0;
    assign data[8329] = 16'b0;
    assign data[8330] = ~16'b0;
    assign data[8331] = ~16'b0;
    assign data[8332] = ~16'b0;
    assign data[8333] = ~16'b0;
    assign data[8334] = ~16'b0;
    assign data[8335] = ~16'b0;
    assign data[8336] = ~16'b0;
    assign data[8337] = ~16'b0;
    assign data[8338] = ~16'b0;
    assign data[8339] = ~16'b0;
    assign data[8340] = ~16'b0;
    assign data[8341] = ~16'b0;
    assign data[8342] = ~16'b0;
    assign data[8343] = ~16'b0;
    assign data[8344] = ~16'b0;
    assign data[8345] = ~16'b0;
    assign data[8346] = ~16'b0;
    assign data[8347] = ~16'b0;
    assign data[8348] = ~16'b0;
    assign data[8349] = ~16'b0;
    assign data[8350] = ~16'b0;
    assign data[8351] = ~16'b0;
    assign data[8352] = ~16'b0;
    assign data[8353] = ~16'b0;
    assign data[8354] = ~16'b0;
    assign data[8355] = ~16'b0;
    assign data[8356] = ~16'b0;
    assign data[8357] = ~16'b0;
    assign data[8358] = ~16'b0;
    assign data[8359] = ~16'b0;
    assign data[8360] = ~16'b0;
    assign data[8361] = ~16'b0;
    assign data[8362] = ~16'b0;
    assign data[8363] = ~16'b0;
    assign data[8364] = ~16'b0;
    assign data[8365] = ~16'b0;
    assign data[8366] = ~16'b0;
    assign data[8367] = ~16'b0;
    assign data[8368] = ~16'b0;
    assign data[8369] = ~16'b0;
    assign data[8370] = ~16'b0;
    assign data[8371] = ~16'b0;
    assign data[8372] = ~16'b0;
    assign data[8373] = ~16'b0;
    assign data[8374] = ~16'b0;
    assign data[8375] = ~16'b0;
    assign data[8376] = ~16'b0;
    assign data[8377] = ~16'b0;
    assign data[8378] = ~16'b0;
    assign data[8379] = ~16'b0;
    assign data[8380] = ~16'b0;
    assign data[8381] = ~16'b0;
    assign data[8382] = ~16'b0;
    assign data[8383] = ~16'b0;
    assign data[8384] = ~16'b0;
    assign data[8385] = ~16'b0;
    assign data[8386] = ~16'b0;
    assign data[8387] = ~16'b0;
    assign data[8388] = ~16'b0;
    assign data[8389] = ~16'b0;
    assign data[8390] = ~16'b0;
    assign data[8391] = ~16'b0;
    assign data[8392] = ~16'b0;
    assign data[8393] = ~16'b0;
    assign data[8394] = ~16'b0;
    assign data[8395] = ~16'b0;
    assign data[8396] = ~16'b0;
    assign data[8397] = ~16'b0;
    assign data[8398] = ~16'b0;
    assign data[8399] = ~16'b0;
    assign data[8400] = ~16'b0;
    assign data[8401] = ~16'b0;
    assign data[8402] = ~16'b0;
    assign data[8403] = ~16'b0;
    assign data[8404] = ~16'b0;
    assign data[8405] = ~16'b0;
    assign data[8406] = ~16'b0;
    assign data[8407] = ~16'b0;
    assign data[8408] = ~16'b0;
    assign data[8409] = ~16'b0;
    assign data[8410] = ~16'b0;
    assign data[8411] = ~16'b0;
    assign data[8412] = ~16'b0;
    assign data[8413] = ~16'b0;
    assign data[8414] = ~16'b0;
    assign data[8415] = ~16'b0;
    assign data[8416] = ~16'b0;
    assign data[8417] = ~16'b0;
    assign data[8418] = ~16'b0;
    assign data[8419] = ~16'b0;
    assign data[8420] = ~16'b0;
    assign data[8421] = ~16'b0;
    assign data[8422] = ~16'b0;
    assign data[8423] = ~16'b0;
    assign data[8424] = ~16'b0;
    assign data[8425] = ~16'b0;
    assign data[8426] = ~16'b0;
    assign data[8427] = ~16'b0;
    assign data[8428] = ~16'b0;
    assign data[8429] = ~16'b0;
    assign data[8430] = ~16'b0;
    assign data[8431] = ~16'b0;
    assign data[8432] = ~16'b0;
    assign data[8433] = ~16'b0;
    assign data[8434] = ~16'b0;
    assign data[8435] = ~16'b0;
    assign data[8436] = ~16'b0;
    assign data[8437] = ~16'b0;
    assign data[8438] = ~16'b0;
    assign data[8439] = ~16'b0;
    assign data[8440] = ~16'b0;
    assign data[8441] = ~16'b0;
    assign data[8442] = ~16'b0;
    assign data[8443] = ~16'b0;
    assign data[8444] = ~16'b0;
    assign data[8445] = ~16'b0;
    assign data[8446] = ~16'b0;
    assign data[8447] = ~16'b0;
    assign data[8448] = ~16'b0;
    assign data[8449] = ~16'b0;
    assign data[8450] = ~16'b0;
    assign data[8451] = ~16'b0;
    assign data[8452] = ~16'b0;
    assign data[8453] = ~16'b0;
    assign data[8454] = ~16'b0;
    assign data[8455] = ~16'b0;
    assign data[8456] = ~16'b0;
    assign data[8457] = ~16'b0;
    assign data[8458] = ~16'b0;
    assign data[8459] = ~16'b0;
    assign data[8460] = ~16'b0;
    assign data[8461] = ~16'b0;
    assign data[8462] = ~16'b0;
    assign data[8463] = ~16'b0;
    assign data[8464] = ~16'b0;
    assign data[8465] = ~16'b0;
    assign data[8466] = ~16'b0;
    assign data[8467] = ~16'b0;
    assign data[8468] = ~16'b0;
    assign data[8469] = ~16'b0;
    assign data[8470] = 16'b0;
    assign data[8471] = 16'b0;
    assign data[8472] = 16'b0;
    assign data[8473] = 16'b0;
    assign data[8474] = 16'b0;
    assign data[8475] = 16'b0;
    assign data[8476] = 16'b0;
    assign data[8477] = 16'b0;
    assign data[8478] = 16'b0;
    assign data[8479] = 16'b0;
    assign data[8480] = 16'b0;
    assign data[8481] = 16'b0;
    assign data[8482] = 16'b0;
    assign data[8483] = 16'b0;
    assign data[8484] = 16'b0;
    assign data[8485] = 16'b0;
    assign data[8486] = 16'b0;
    assign data[8487] = 16'b0;
    assign data[8488] = 16'b0;
    assign data[8489] = 16'b0;
    assign data[8490] = 16'b0;
    assign data[8491] = 16'b0;
    assign data[8492] = ~16'b0;
    assign data[8493] = ~16'b0;
    assign data[8494] = ~16'b0;
    assign data[8495] = ~16'b0;
    assign data[8496] = ~16'b0;
    assign data[8497] = ~16'b0;
    assign data[8498] = ~16'b0;
    assign data[8499] = ~16'b0;
    assign data[8500] = 16'b0;
    assign data[8501] = 16'b0;
    assign data[8502] = ~16'b0;
    assign data[8503] = ~16'b0;
    assign data[8504] = ~16'b0;
    assign data[8505] = ~16'b0;
    assign data[8506] = ~16'b0;
    assign data[8507] = ~16'b0;
    assign data[8508] = ~16'b0;
    assign data[8509] = ~16'b0;
    assign data[8510] = 16'b0;
    assign data[8511] = 16'b0;
    assign data[8512] = ~16'b0;
    assign data[8513] = ~16'b0;
    assign data[8514] = ~16'b0;
    assign data[8515] = ~16'b0;
    assign data[8516] = ~16'b0;
    assign data[8517] = ~16'b0;
    assign data[8518] = ~16'b0;
    assign data[8519] = ~16'b0;
    assign data[8520] = 16'b0;
    assign data[8521] = 16'b0;
    assign data[8522] = ~16'b0;
    assign data[8523] = ~16'b0;
    assign data[8524] = ~16'b0;
    assign data[8525] = ~16'b0;
    assign data[8526] = ~16'b0;
    assign data[8527] = ~16'b0;
    assign data[8528] = ~16'b0;
    assign data[8529] = ~16'b0;
    assign data[8530] = 16'b0;
    assign data[8531] = 16'b0;
    assign data[8532] = ~16'b0;
    assign data[8533] = ~16'b0;
    assign data[8534] = ~16'b0;
    assign data[8535] = ~16'b0;
    assign data[8536] = ~16'b0;
    assign data[8537] = ~16'b0;
    assign data[8538] = ~16'b0;
    assign data[8539] = ~16'b0;
    assign data[8540] = 16'b0;
    assign data[8541] = 16'b0;
    assign data[8542] = ~16'b0;
    assign data[8543] = ~16'b0;
    assign data[8544] = ~16'b0;
    assign data[8545] = ~16'b0;
    assign data[8546] = ~16'b0;
    assign data[8547] = ~16'b0;
    assign data[8548] = ~16'b0;
    assign data[8549] = ~16'b0;
    assign data[8550] = 16'b0;
    assign data[8551] = 16'b0;
    assign data[8552] = ~16'b0;
    assign data[8553] = ~16'b0;
    assign data[8554] = ~16'b0;
    assign data[8555] = ~16'b0;
    assign data[8556] = ~16'b0;
    assign data[8557] = ~16'b0;
    assign data[8558] = ~16'b0;
    assign data[8559] = ~16'b0;
    assign data[8560] = 16'b0;
    assign data[8561] = 16'b0;
    assign data[8562] = ~16'b0;
    assign data[8563] = ~16'b0;
    assign data[8564] = ~16'b0;
    assign data[8565] = ~16'b0;
    assign data[8566] = ~16'b0;
    assign data[8567] = ~16'b0;
    assign data[8568] = ~16'b0;
    assign data[8569] = ~16'b0;
    assign data[8570] = 16'b0;
    assign data[8571] = 16'b0;
    assign data[8572] = ~16'b0;
    assign data[8573] = ~16'b0;
    assign data[8574] = ~16'b0;
    assign data[8575] = ~16'b0;
    assign data[8576] = ~16'b0;
    assign data[8577] = ~16'b0;
    assign data[8578] = ~16'b0;
    assign data[8579] = ~16'b0;
    assign data[8580] = 16'b0;
    assign data[8581] = 16'b0;
    assign data[8582] = ~16'b0;
    assign data[8583] = ~16'b0;
    assign data[8584] = ~16'b0;
    assign data[8585] = ~16'b0;
    assign data[8586] = ~16'b0;
    assign data[8587] = ~16'b0;
    assign data[8588] = ~16'b0;
    assign data[8589] = ~16'b0;
    assign data[8590] = 16'b0;
    assign data[8591] = 16'b0;
    assign data[8592] = ~16'b0;
    assign data[8593] = ~16'b0;
    assign data[8594] = ~16'b0;
    assign data[8595] = ~16'b0;
    assign data[8596] = ~16'b0;
    assign data[8597] = ~16'b0;
    assign data[8598] = ~16'b0;
    assign data[8599] = ~16'b0;
    assign data[8600] = 16'b0;
    assign data[8601] = 16'b0;
    assign data[8602] = ~16'b0;
    assign data[8603] = ~16'b0;
    assign data[8604] = ~16'b0;
    assign data[8605] = ~16'b0;
    assign data[8606] = ~16'b0;
    assign data[8607] = ~16'b0;
    assign data[8608] = ~16'b0;
    assign data[8609] = ~16'b0;
    assign data[8610] = 16'b0;
    assign data[8611] = 16'b0;
    assign data[8612] = ~16'b0;
    assign data[8613] = ~16'b0;
    assign data[8614] = ~16'b0;
    assign data[8615] = ~16'b0;
    assign data[8616] = ~16'b0;
    assign data[8617] = ~16'b0;
    assign data[8618] = ~16'b0;
    assign data[8619] = ~16'b0;
    assign data[8620] = 16'b0;
    assign data[8621] = 16'b0;
    assign data[8622] = ~16'b0;
    assign data[8623] = ~16'b0;
    assign data[8624] = ~16'b0;
    assign data[8625] = ~16'b0;
    assign data[8626] = ~16'b0;
    assign data[8627] = ~16'b0;
    assign data[8628] = ~16'b0;
    assign data[8629] = ~16'b0;
    assign data[8630] = 16'b0;
    assign data[8631] = 16'b0;
    assign data[8632] = ~16'b0;
    assign data[8633] = ~16'b0;
    assign data[8634] = ~16'b0;
    assign data[8635] = ~16'b0;
    assign data[8636] = ~16'b0;
    assign data[8637] = ~16'b0;
    assign data[8638] = ~16'b0;
    assign data[8639] = ~16'b0;
    assign data[8640] = 16'b0;
    assign data[8641] = 16'b0;
    assign data[8642] = ~16'b0;
    assign data[8643] = ~16'b0;
    assign data[8644] = ~16'b0;
    assign data[8645] = ~16'b0;
    assign data[8646] = ~16'b0;
    assign data[8647] = ~16'b0;
    assign data[8648] = ~16'b0;
    assign data[8649] = ~16'b0;
    assign data[8650] = 16'b0;
    assign data[8651] = 16'b0;
    assign data[8652] = ~16'b0;
    assign data[8653] = ~16'b0;
    assign data[8654] = ~16'b0;
    assign data[8655] = ~16'b0;
    assign data[8656] = ~16'b0;
    assign data[8657] = ~16'b0;
    assign data[8658] = ~16'b0;
    assign data[8659] = ~16'b0;
    assign data[8660] = 16'b0;
    assign data[8661] = 16'b0;
    assign data[8662] = ~16'b0;
    assign data[8663] = ~16'b0;
    assign data[8664] = ~16'b0;
    assign data[8665] = ~16'b0;
    assign data[8666] = ~16'b0;
    assign data[8667] = ~16'b0;
    assign data[8668] = ~16'b0;
    assign data[8669] = ~16'b0;
    assign data[8670] = 16'b0;
    assign data[8671] = 16'b0;
    assign data[8672] = ~16'b0;
    assign data[8673] = ~16'b0;
    assign data[8674] = ~16'b0;
    assign data[8675] = ~16'b0;
    assign data[8676] = ~16'b0;
    assign data[8677] = ~16'b0;
    assign data[8678] = ~16'b0;
    assign data[8679] = ~16'b0;
    assign data[8680] = 16'b0;
    assign data[8681] = 16'b0;
    assign data[8682] = ~16'b0;
    assign data[8683] = ~16'b0;
    assign data[8684] = ~16'b0;
    assign data[8685] = ~16'b0;
    assign data[8686] = ~16'b0;
    assign data[8687] = ~16'b0;
    assign data[8688] = ~16'b0;
    assign data[8689] = ~16'b0;
    assign data[8690] = 16'b0;
    assign data[8691] = 16'b0;
    assign data[8692] = 16'b0;
    assign data[8693] = 16'b0;
    assign data[8694] = 16'b0;
    assign data[8695] = 16'b0;
    assign data[8696] = 16'b0;
    assign data[8697] = 16'b0;
    assign data[8698] = 16'b0;
    assign data[8699] = 16'b0;
    assign data[8700] = 16'b0;
    assign data[8701] = 16'b0;
    assign data[8702] = 16'b0;
    assign data[8703] = 16'b0;
    assign data[8704] = 16'b0;
    assign data[8705] = 16'b0;
    assign data[8706] = 16'b0;
    assign data[8707] = 16'b0;
    assign data[8708] = 16'b0;
    assign data[8709] = 16'b0;
    assign data[8710] = ~16'b0;
    assign data[8711] = ~16'b0;
    assign data[8712] = ~16'b0;
    assign data[8713] = ~16'b0;
    assign data[8714] = ~16'b0;
    assign data[8715] = ~16'b0;
    assign data[8716] = ~16'b0;
    assign data[8717] = ~16'b0;
    assign data[8718] = ~16'b0;
    assign data[8719] = ~16'b0;
    assign data[8720] = ~16'b0;
    assign data[8721] = ~16'b0;
    assign data[8722] = ~16'b0;
    assign data[8723] = ~16'b0;
    assign data[8724] = ~16'b0;
    assign data[8725] = ~16'b0;
    assign data[8726] = ~16'b0;
    assign data[8727] = ~16'b0;
    assign data[8728] = ~16'b0;
    assign data[8729] = ~16'b0;
    assign data[8730] = ~16'b0;
    assign data[8731] = ~16'b0;
    assign data[8732] = ~16'b0;
    assign data[8733] = ~16'b0;
    assign data[8734] = ~16'b0;
    assign data[8735] = ~16'b0;
    assign data[8736] = ~16'b0;
    assign data[8737] = ~16'b0;
    assign data[8738] = ~16'b0;
    assign data[8739] = ~16'b0;
    assign data[8740] = ~16'b0;
    assign data[8741] = ~16'b0;
    assign data[8742] = ~16'b0;
    assign data[8743] = ~16'b0;
    assign data[8744] = ~16'b0;
    assign data[8745] = ~16'b0;
    assign data[8746] = ~16'b0;
    assign data[8747] = ~16'b0;
    assign data[8748] = ~16'b0;
    assign data[8749] = ~16'b0;
    assign data[8750] = ~16'b0;
    assign data[8751] = ~16'b0;
    assign data[8752] = ~16'b0;
    assign data[8753] = ~16'b0;
    assign data[8754] = ~16'b0;
    assign data[8755] = ~16'b0;
    assign data[8756] = ~16'b0;
    assign data[8757] = ~16'b0;
    assign data[8758] = ~16'b0;
    assign data[8759] = ~16'b0;
    assign data[8760] = ~16'b0;
    assign data[8761] = ~16'b0;
    assign data[8762] = ~16'b0;
    assign data[8763] = ~16'b0;
    assign data[8764] = ~16'b0;
    assign data[8765] = ~16'b0;
    assign data[8766] = ~16'b0;
    assign data[8767] = ~16'b0;
    assign data[8768] = ~16'b0;
    assign data[8769] = ~16'b0;
    assign data[8770] = ~16'b0;
    assign data[8771] = ~16'b0;
    assign data[8772] = ~16'b0;
    assign data[8773] = ~16'b0;
    assign data[8774] = ~16'b0;
    assign data[8775] = ~16'b0;
    assign data[8776] = ~16'b0;
    assign data[8777] = ~16'b0;
    assign data[8778] = ~16'b0;
    assign data[8779] = ~16'b0;
    assign data[8780] = ~16'b0;
    assign data[8781] = ~16'b0;
    assign data[8782] = ~16'b0;
    assign data[8783] = ~16'b0;
    assign data[8784] = ~16'b0;
    assign data[8785] = ~16'b0;
    assign data[8786] = ~16'b0;
    assign data[8787] = ~16'b0;
    assign data[8788] = ~16'b0;
    assign data[8789] = ~16'b0;
    assign data[8790] = ~16'b0;
    assign data[8791] = ~16'b0;
    assign data[8792] = ~16'b0;
    assign data[8793] = ~16'b0;
    assign data[8794] = ~16'b0;
    assign data[8795] = ~16'b0;
    assign data[8796] = ~16'b0;
    assign data[8797] = ~16'b0;
    assign data[8798] = ~16'b0;
    assign data[8799] = ~16'b0;
    assign data[8800] = ~16'b0;
    assign data[8801] = ~16'b0;
    assign data[8802] = ~16'b0;
    assign data[8803] = ~16'b0;
    assign data[8804] = ~16'b0;
    assign data[8805] = ~16'b0;
    assign data[8806] = ~16'b0;
    assign data[8807] = ~16'b0;
    assign data[8808] = ~16'b0;
    assign data[8809] = ~16'b0;
    assign data[8810] = ~16'b0;
    assign data[8811] = ~16'b0;
    assign data[8812] = ~16'b0;
    assign data[8813] = ~16'b0;
    assign data[8814] = ~16'b0;
    assign data[8815] = ~16'b0;
    assign data[8816] = ~16'b0;
    assign data[8817] = ~16'b0;
    assign data[8818] = ~16'b0;
    assign data[8819] = ~16'b0;
    assign data[8820] = ~16'b0;
    assign data[8821] = ~16'b0;
    assign data[8822] = ~16'b0;
    assign data[8823] = ~16'b0;
    assign data[8824] = ~16'b0;
    assign data[8825] = ~16'b0;
    assign data[8826] = ~16'b0;
    assign data[8827] = ~16'b0;
    assign data[8828] = ~16'b0;
    assign data[8829] = ~16'b0;
    assign data[8830] = ~16'b0;
    assign data[8831] = ~16'b0;
    assign data[8832] = ~16'b0;
    assign data[8833] = ~16'b0;
    assign data[8834] = ~16'b0;
    assign data[8835] = ~16'b0;
    assign data[8836] = ~16'b0;
    assign data[8837] = ~16'b0;
    assign data[8838] = ~16'b0;
    assign data[8839] = ~16'b0;
    assign data[8840] = ~16'b0;
    assign data[8841] = ~16'b0;
    assign data[8842] = ~16'b0;
    assign data[8843] = ~16'b0;
    assign data[8844] = ~16'b0;
    assign data[8845] = ~16'b0;
    assign data[8846] = ~16'b0;
    assign data[8847] = ~16'b0;
    assign data[8848] = ~16'b0;
    assign data[8849] = ~16'b0;
    assign data[8850] = ~16'b0;
    assign data[8851] = ~16'b0;
    assign data[8852] = ~16'b0;
    assign data[8853] = ~16'b0;
    assign data[8854] = ~16'b0;
    assign data[8855] = ~16'b0;
    assign data[8856] = ~16'b0;
    assign data[8857] = ~16'b0;
    assign data[8858] = ~16'b0;
    assign data[8859] = ~16'b0;
    assign data[8860] = 16'b0;
    assign data[8861] = 16'b0;
    assign data[8862] = 16'b0;
    assign data[8863] = 16'b0;
    assign data[8864] = 16'b0;
    assign data[8865] = 16'b0;
    assign data[8866] = 16'b0;
    assign data[8867] = 16'b0;
    assign data[8868] = 16'b0;
    assign data[8869] = 16'b0;
    assign data[8870] = 16'b0;
    assign data[8871] = 16'b0;
    assign data[8872] = 16'b0;
    assign data[8873] = 16'b0;
    assign data[8874] = 16'b0;
    assign data[8875] = 16'b0;
    assign data[8876] = 16'b0;
    assign data[8877] = 16'b0;
    assign data[8878] = 16'b0;
    assign data[8879] = 16'b0;
    assign data[8880] = 16'b0;
    assign data[8881] = 16'b0;
    assign data[8882] = ~16'b0;
    assign data[8883] = ~16'b0;
    assign data[8884] = ~16'b0;
    assign data[8885] = ~16'b0;
    assign data[8886] = ~16'b0;
    assign data[8887] = ~16'b0;
    assign data[8888] = ~16'b0;
    assign data[8889] = ~16'b0;
    assign data[8890] = 16'b0;
    assign data[8891] = 16'b0;
    assign data[8892] = ~16'b0;
    assign data[8893] = ~16'b0;
    assign data[8894] = ~16'b0;
    assign data[8895] = ~16'b0;
    assign data[8896] = ~16'b0;
    assign data[8897] = ~16'b0;
    assign data[8898] = ~16'b0;
    assign data[8899] = ~16'b0;
    assign data[8900] = 16'b0;
    assign data[8901] = 16'b0;
    assign data[8902] = ~16'b0;
    assign data[8903] = ~16'b0;
    assign data[8904] = ~16'b0;
    assign data[8905] = ~16'b0;
    assign data[8906] = ~16'b0;
    assign data[8907] = ~16'b0;
    assign data[8908] = ~16'b0;
    assign data[8909] = ~16'b0;
    assign data[8910] = 16'b0;
    assign data[8911] = 16'b0;
    assign data[8912] = ~16'b0;
    assign data[8913] = ~16'b0;
    assign data[8914] = ~16'b0;
    assign data[8915] = ~16'b0;
    assign data[8916] = ~16'b0;
    assign data[8917] = ~16'b0;
    assign data[8918] = ~16'b0;
    assign data[8919] = ~16'b0;
    assign data[8920] = 16'b0;
    assign data[8921] = 16'b0;
    assign data[8922] = ~16'b0;
    assign data[8923] = ~16'b0;
    assign data[8924] = ~16'b0;
    assign data[8925] = ~16'b0;
    assign data[8926] = ~16'b0;
    assign data[8927] = ~16'b0;
    assign data[8928] = ~16'b0;
    assign data[8929] = ~16'b0;
    assign data[8930] = 16'b0;
    assign data[8931] = 16'b0;
    assign data[8932] = ~16'b0;
    assign data[8933] = ~16'b0;
    assign data[8934] = ~16'b0;
    assign data[8935] = ~16'b0;
    assign data[8936] = ~16'b0;
    assign data[8937] = ~16'b0;
    assign data[8938] = ~16'b0;
    assign data[8939] = ~16'b0;
    assign data[8940] = 16'b0;
    assign data[8941] = 16'b0;
    assign data[8942] = ~16'b0;
    assign data[8943] = ~16'b0;
    assign data[8944] = ~16'b0;
    assign data[8945] = ~16'b0;
    assign data[8946] = ~16'b0;
    assign data[8947] = ~16'b0;
    assign data[8948] = ~16'b0;
    assign data[8949] = ~16'b0;
    assign data[8950] = 16'b0;
    assign data[8951] = 16'b0;
    assign data[8952] = ~16'b0;
    assign data[8953] = ~16'b0;
    assign data[8954] = ~16'b0;
    assign data[8955] = ~16'b0;
    assign data[8956] = ~16'b0;
    assign data[8957] = ~16'b0;
    assign data[8958] = ~16'b0;
    assign data[8959] = ~16'b0;
    assign data[8960] = 16'b0;
    assign data[8961] = 16'b0;
    assign data[8962] = ~16'b0;
    assign data[8963] = ~16'b0;
    assign data[8964] = ~16'b0;
    assign data[8965] = ~16'b0;
    assign data[8966] = ~16'b0;
    assign data[8967] = ~16'b0;
    assign data[8968] = ~16'b0;
    assign data[8969] = ~16'b0;
    assign data[8970] = 16'b0;
    assign data[8971] = 16'b0;
    assign data[8972] = ~16'b0;
    assign data[8973] = ~16'b0;
    assign data[8974] = ~16'b0;
    assign data[8975] = ~16'b0;
    assign data[8976] = ~16'b0;
    assign data[8977] = ~16'b0;
    assign data[8978] = ~16'b0;
    assign data[8979] = ~16'b0;
    assign data[8980] = 16'b0;
    assign data[8981] = 16'b0;
    assign data[8982] = ~16'b0;
    assign data[8983] = ~16'b0;
    assign data[8984] = ~16'b0;
    assign data[8985] = ~16'b0;
    assign data[8986] = ~16'b0;
    assign data[8987] = ~16'b0;
    assign data[8988] = ~16'b0;
    assign data[8989] = ~16'b0;
    assign data[8990] = 16'b0;
    assign data[8991] = 16'b0;
    assign data[8992] = ~16'b0;
    assign data[8993] = ~16'b0;
    assign data[8994] = ~16'b0;
    assign data[8995] = ~16'b0;
    assign data[8996] = ~16'b0;
    assign data[8997] = ~16'b0;
    assign data[8998] = ~16'b0;
    assign data[8999] = ~16'b0;
    assign data[9000] = 16'b0;
    assign data[9001] = 16'b0;
    assign data[9002] = ~16'b0;
    assign data[9003] = ~16'b0;
    assign data[9004] = ~16'b0;
    assign data[9005] = ~16'b0;
    assign data[9006] = ~16'b0;
    assign data[9007] = ~16'b0;
    assign data[9008] = ~16'b0;
    assign data[9009] = ~16'b0;
    assign data[9010] = 16'b0;
    assign data[9011] = 16'b0;
    assign data[9012] = ~16'b0;
    assign data[9013] = ~16'b0;
    assign data[9014] = ~16'b0;
    assign data[9015] = ~16'b0;
    assign data[9016] = ~16'b0;
    assign data[9017] = ~16'b0;
    assign data[9018] = ~16'b0;
    assign data[9019] = ~16'b0;
    assign data[9020] = 16'b0;
    assign data[9021] = 16'b0;
    assign data[9022] = ~16'b0;
    assign data[9023] = ~16'b0;
    assign data[9024] = ~16'b0;
    assign data[9025] = ~16'b0;
    assign data[9026] = ~16'b0;
    assign data[9027] = ~16'b0;
    assign data[9028] = ~16'b0;
    assign data[9029] = ~16'b0;
    assign data[9030] = 16'b0;
    assign data[9031] = 16'b0;
    assign data[9032] = ~16'b0;
    assign data[9033] = ~16'b0;
    assign data[9034] = ~16'b0;
    assign data[9035] = ~16'b0;
    assign data[9036] = ~16'b0;
    assign data[9037] = ~16'b0;
    assign data[9038] = ~16'b0;
    assign data[9039] = ~16'b0;
    assign data[9040] = 16'b0;
    assign data[9041] = 16'b0;
    assign data[9042] = ~16'b0;
    assign data[9043] = ~16'b0;
    assign data[9044] = ~16'b0;
    assign data[9045] = ~16'b0;
    assign data[9046] = ~16'b0;
    assign data[9047] = ~16'b0;
    assign data[9048] = ~16'b0;
    assign data[9049] = ~16'b0;
    assign data[9050] = 16'b0;
    assign data[9051] = 16'b0;
    assign data[9052] = ~16'b0;
    assign data[9053] = ~16'b0;
    assign data[9054] = ~16'b0;
    assign data[9055] = ~16'b0;
    assign data[9056] = ~16'b0;
    assign data[9057] = ~16'b0;
    assign data[9058] = ~16'b0;
    assign data[9059] = ~16'b0;
    assign data[9060] = 16'b0;
    assign data[9061] = 16'b0;
    assign data[9062] = ~16'b0;
    assign data[9063] = ~16'b0;
    assign data[9064] = ~16'b0;
    assign data[9065] = ~16'b0;
    assign data[9066] = ~16'b0;
    assign data[9067] = ~16'b0;
    assign data[9068] = ~16'b0;
    assign data[9069] = ~16'b0;
    assign data[9070] = 16'b0;
    assign data[9071] = 16'b0;
    assign data[9072] = ~16'b0;
    assign data[9073] = ~16'b0;
    assign data[9074] = ~16'b0;
    assign data[9075] = ~16'b0;
    assign data[9076] = ~16'b0;
    assign data[9077] = ~16'b0;
    assign data[9078] = ~16'b0;
    assign data[9079] = ~16'b0;
    assign data[9080] = 16'b0;
    assign data[9081] = 16'b0;
    assign data[9082] = ~16'b0;
    assign data[9083] = ~16'b0;
    assign data[9084] = ~16'b0;
    assign data[9085] = ~16'b0;
    assign data[9086] = ~16'b0;
    assign data[9087] = ~16'b0;
    assign data[9088] = ~16'b0;
    assign data[9089] = ~16'b0;
    assign data[9090] = 16'b0;
    assign data[9091] = 16'b0;
    assign data[9092] = ~16'b0;
    assign data[9093] = ~16'b0;
    assign data[9094] = ~16'b0;
    assign data[9095] = ~16'b0;
    assign data[9096] = ~16'b0;
    assign data[9097] = ~16'b0;
    assign data[9098] = ~16'b0;
    assign data[9099] = ~16'b0;
    assign data[9100] = 16'b0;
    assign data[9101] = 16'b0;
    assign data[9102] = ~16'b0;
    assign data[9103] = ~16'b0;
    assign data[9104] = ~16'b0;
    assign data[9105] = ~16'b0;
    assign data[9106] = ~16'b0;
    assign data[9107] = ~16'b0;
    assign data[9108] = ~16'b0;
    assign data[9109] = ~16'b0;
    assign data[9110] = 16'b0;
    assign data[9111] = 16'b0;
    assign data[9112] = ~16'b0;
    assign data[9113] = ~16'b0;
    assign data[9114] = ~16'b0;
    assign data[9115] = ~16'b0;
    assign data[9116] = ~16'b0;
    assign data[9117] = ~16'b0;
    assign data[9118] = ~16'b0;
    assign data[9119] = ~16'b0;
    assign data[9120] = 16'b0;
    assign data[9121] = 16'b0;
    assign data[9122] = ~16'b0;
    assign data[9123] = ~16'b0;
    assign data[9124] = ~16'b0;
    assign data[9125] = ~16'b0;
    assign data[9126] = ~16'b0;
    assign data[9127] = ~16'b0;
    assign data[9128] = ~16'b0;
    assign data[9129] = ~16'b0;
    assign data[9130] = 16'b0;
    assign data[9131] = 16'b0;
    assign data[9132] = ~16'b0;
    assign data[9133] = ~16'b0;
    assign data[9134] = ~16'b0;
    assign data[9135] = ~16'b0;
    assign data[9136] = ~16'b0;
    assign data[9137] = ~16'b0;
    assign data[9138] = ~16'b0;
    assign data[9139] = ~16'b0;
    assign data[9140] = 16'b0;
    assign data[9141] = 16'b0;
    assign data[9142] = ~16'b0;
    assign data[9143] = ~16'b0;
    assign data[9144] = ~16'b0;
    assign data[9145] = ~16'b0;
    assign data[9146] = ~16'b0;
    assign data[9147] = ~16'b0;
    assign data[9148] = ~16'b0;
    assign data[9149] = ~16'b0;
    assign data[9150] = 16'b0;
    assign data[9151] = 16'b0;
    assign data[9152] = ~16'b0;
    assign data[9153] = ~16'b0;
    assign data[9154] = ~16'b0;
    assign data[9155] = ~16'b0;
    assign data[9156] = ~16'b0;
    assign data[9157] = ~16'b0;
    assign data[9158] = ~16'b0;
    assign data[9159] = ~16'b0;
    assign data[9160] = 16'b0;
    assign data[9161] = 16'b0;
    assign data[9162] = ~16'b0;
    assign data[9163] = ~16'b0;
    assign data[9164] = ~16'b0;
    assign data[9165] = ~16'b0;
    assign data[9166] = ~16'b0;
    assign data[9167] = ~16'b0;
    assign data[9168] = ~16'b0;
    assign data[9169] = ~16'b0;
    assign data[9170] = 16'b0;
    assign data[9171] = 16'b0;
    assign data[9172] = ~16'b0;
    assign data[9173] = ~16'b0;
    assign data[9174] = ~16'b0;
    assign data[9175] = ~16'b0;
    assign data[9176] = ~16'b0;
    assign data[9177] = ~16'b0;
    assign data[9178] = ~16'b0;
    assign data[9179] = ~16'b0;
    assign data[9180] = 16'b0;
    assign data[9181] = 16'b0;
    assign data[9182] = ~16'b0;
    assign data[9183] = ~16'b0;
    assign data[9184] = ~16'b0;
    assign data[9185] = ~16'b0;
    assign data[9186] = ~16'b0;
    assign data[9187] = ~16'b0;
    assign data[9188] = ~16'b0;
    assign data[9189] = ~16'b0;
    assign data[9190] = 16'b0;
    assign data[9191] = 16'b0;
    assign data[9192] = ~16'b0;
    assign data[9193] = ~16'b0;
    assign data[9194] = ~16'b0;
    assign data[9195] = ~16'b0;
    assign data[9196] = ~16'b0;
    assign data[9197] = ~16'b0;
    assign data[9198] = ~16'b0;
    assign data[9199] = ~16'b0;
    assign data[9200] = 16'b0;
    assign data[9201] = 16'b0;
    assign data[9202] = ~16'b0;
    assign data[9203] = ~16'b0;
    assign data[9204] = ~16'b0;
    assign data[9205] = ~16'b0;
    assign data[9206] = ~16'b0;
    assign data[9207] = ~16'b0;
    assign data[9208] = ~16'b0;
    assign data[9209] = ~16'b0;
    assign data[9210] = 16'b0;
    assign data[9211] = 16'b0;
    assign data[9212] = ~16'b0;
    assign data[9213] = ~16'b0;
    assign data[9214] = ~16'b0;
    assign data[9215] = ~16'b0;
    assign data[9216] = ~16'b0;
    assign data[9217] = ~16'b0;
    assign data[9218] = ~16'b0;
    assign data[9219] = ~16'b0;
    assign data[9220] = 16'b0;
    assign data[9221] = 16'b0;
    assign data[9222] = 16'b0;
    assign data[9223] = 16'b0;
    assign data[9224] = 16'b0;
    assign data[9225] = 16'b0;
    assign data[9226] = 16'b0;
    assign data[9227] = 16'b0;
    assign data[9228] = 16'b0;
    assign data[9229] = 16'b0;
    assign data[9230] = 16'b0;
    assign data[9231] = 16'b0;
    assign data[9232] = 16'b0;
    assign data[9233] = 16'b0;
    assign data[9234] = 16'b0;
    assign data[9235] = 16'b0;
    assign data[9236] = 16'b0;
    assign data[9237] = 16'b0;
    assign data[9238] = 16'b0;
    assign data[9239] = 16'b0;
    assign data[9240] = ~16'b0;
    assign data[9241] = ~16'b0;
    assign data[9242] = ~16'b0;
    assign data[9243] = ~16'b0;
    assign data[9244] = ~16'b0;
    assign data[9245] = ~16'b0;
    assign data[9246] = ~16'b0;
    assign data[9247] = ~16'b0;
    assign data[9248] = ~16'b0;
    assign data[9249] = ~16'b0;
    assign data[9250] = ~16'b0;
    assign data[9251] = ~16'b0;
    assign data[9252] = ~16'b0;
    assign data[9253] = ~16'b0;
    assign data[9254] = ~16'b0;
    assign data[9255] = ~16'b0;
    assign data[9256] = ~16'b0;
    assign data[9257] = ~16'b0;
    assign data[9258] = ~16'b0;
    assign data[9259] = ~16'b0;
    assign data[9260] = ~16'b0;
    assign data[9261] = ~16'b0;
    assign data[9262] = ~16'b0;
    assign data[9263] = ~16'b0;
    assign data[9264] = ~16'b0;
    assign data[9265] = ~16'b0;
    assign data[9266] = ~16'b0;
    assign data[9267] = ~16'b0;
    assign data[9268] = ~16'b0;
    assign data[9269] = ~16'b0;
    assign data[9270] = ~16'b0;
    assign data[9271] = ~16'b0;
    assign data[9272] = ~16'b0;
    assign data[9273] = ~16'b0;
    assign data[9274] = ~16'b0;
    assign data[9275] = ~16'b0;
    assign data[9276] = ~16'b0;
    assign data[9277] = ~16'b0;
    assign data[9278] = ~16'b0;
    assign data[9279] = ~16'b0;
    assign data[9280] = ~16'b0;
    assign data[9281] = ~16'b0;
    assign data[9282] = ~16'b0;
    assign data[9283] = ~16'b0;
    assign data[9284] = ~16'b0;
    assign data[9285] = ~16'b0;
    assign data[9286] = ~16'b0;
    assign data[9287] = ~16'b0;
    assign data[9288] = ~16'b0;
    assign data[9289] = ~16'b0;
    assign data[9290] = ~16'b0;
    assign data[9291] = ~16'b0;
    assign data[9292] = ~16'b0;
    assign data[9293] = ~16'b0;
    assign data[9294] = ~16'b0;
    assign data[9295] = ~16'b0;
    assign data[9296] = ~16'b0;
    assign data[9297] = ~16'b0;
    assign data[9298] = ~16'b0;
    assign data[9299] = ~16'b0;
    assign data[9300] = ~16'b0;
    assign data[9301] = ~16'b0;
    assign data[9302] = ~16'b0;
    assign data[9303] = ~16'b0;
    assign data[9304] = ~16'b0;
    assign data[9305] = ~16'b0;
    assign data[9306] = ~16'b0;
    assign data[9307] = ~16'b0;
    assign data[9308] = ~16'b0;
    assign data[9309] = ~16'b0;
    assign data[9310] = ~16'b0;
    assign data[9311] = ~16'b0;
    assign data[9312] = ~16'b0;
    assign data[9313] = ~16'b0;
    assign data[9314] = ~16'b0;
    assign data[9315] = ~16'b0;
    assign data[9316] = ~16'b0;
    assign data[9317] = ~16'b0;
    assign data[9318] = ~16'b0;
    assign data[9319] = ~16'b0;
    assign data[9320] = ~16'b0;
    assign data[9321] = ~16'b0;
    assign data[9322] = ~16'b0;
    assign data[9323] = ~16'b0;
    assign data[9324] = ~16'b0;
    assign data[9325] = ~16'b0;
    assign data[9326] = ~16'b0;
    assign data[9327] = ~16'b0;
    assign data[9328] = ~16'b0;
    assign data[9329] = ~16'b0;
    assign data[9330] = ~16'b0;
    assign data[9331] = ~16'b0;
    assign data[9332] = ~16'b0;
    assign data[9333] = ~16'b0;
    assign data[9334] = ~16'b0;
    assign data[9335] = ~16'b0;
    assign data[9336] = ~16'b0;
    assign data[9337] = ~16'b0;
    assign data[9338] = ~16'b0;
    assign data[9339] = ~16'b0;
    assign data[9340] = ~16'b0;
    assign data[9341] = ~16'b0;
    assign data[9342] = ~16'b0;
    assign data[9343] = ~16'b0;
    assign data[9344] = ~16'b0;
    assign data[9345] = ~16'b0;
    assign data[9346] = ~16'b0;
    assign data[9347] = ~16'b0;
    assign data[9348] = ~16'b0;
    assign data[9349] = ~16'b0;
    assign data[9350] = ~16'b0;
    assign data[9351] = ~16'b0;
    assign data[9352] = ~16'b0;
    assign data[9353] = ~16'b0;
    assign data[9354] = ~16'b0;
    assign data[9355] = ~16'b0;
    assign data[9356] = ~16'b0;
    assign data[9357] = ~16'b0;
    assign data[9358] = ~16'b0;
    assign data[9359] = ~16'b0;
    assign data[9360] = ~16'b0;
    assign data[9361] = ~16'b0;
    assign data[9362] = ~16'b0;
    assign data[9363] = ~16'b0;
    assign data[9364] = ~16'b0;
    assign data[9365] = ~16'b0;
    assign data[9366] = ~16'b0;
    assign data[9367] = ~16'b0;
    assign data[9368] = ~16'b0;
    assign data[9369] = ~16'b0;
    assign data[9370] = ~16'b0;
    assign data[9371] = ~16'b0;
    assign data[9372] = ~16'b0;
    assign data[9373] = ~16'b0;
    assign data[9374] = ~16'b0;
    assign data[9375] = ~16'b0;
    assign data[9376] = ~16'b0;
    assign data[9377] = ~16'b0;
    assign data[9378] = ~16'b0;
    assign data[9379] = ~16'b0;
    assign data[9380] = ~16'b0;
    assign data[9381] = ~16'b0;
    assign data[9382] = ~16'b0;
    assign data[9383] = ~16'b0;
    assign data[9384] = ~16'b0;
    assign data[9385] = ~16'b0;
    assign data[9386] = ~16'b0;
    assign data[9387] = ~16'b0;
    assign data[9388] = ~16'b0;
    assign data[9389] = ~16'b0;
    assign data[9390] = ~16'b0;
    assign data[9391] = ~16'b0;
    assign data[9392] = ~16'b0;
    assign data[9393] = ~16'b0;
    assign data[9394] = ~16'b0;
    assign data[9395] = ~16'b0;
    assign data[9396] = ~16'b0;
    assign data[9397] = ~16'b0;
    assign data[9398] = ~16'b0;
    assign data[9399] = ~16'b0;
    assign data[9400] = ~16'b0;
    assign data[9401] = ~16'b0;
    assign data[9402] = ~16'b0;
    assign data[9403] = ~16'b0;
    assign data[9404] = ~16'b0;
    assign data[9405] = ~16'b0;
    assign data[9406] = ~16'b0;
    assign data[9407] = ~16'b0;
    assign data[9408] = ~16'b0;
    assign data[9409] = ~16'b0;
    assign data[9410] = ~16'b0;
    assign data[9411] = ~16'b0;
    assign data[9412] = ~16'b0;
    assign data[9413] = ~16'b0;
    assign data[9414] = ~16'b0;
    assign data[9415] = ~16'b0;
    assign data[9416] = ~16'b0;
    assign data[9417] = ~16'b0;
    assign data[9418] = ~16'b0;
    assign data[9419] = ~16'b0;
    assign data[9420] = ~16'b0;
    assign data[9421] = ~16'b0;
    assign data[9422] = ~16'b0;
    assign data[9423] = ~16'b0;
    assign data[9424] = ~16'b0;
    assign data[9425] = ~16'b0;
    assign data[9426] = ~16'b0;
    assign data[9427] = ~16'b0;
    assign data[9428] = ~16'b0;
    assign data[9429] = ~16'b0;
    assign data[9430] = ~16'b0;
    assign data[9431] = ~16'b0;
    assign data[9432] = ~16'b0;
    assign data[9433] = ~16'b0;
    assign data[9434] = ~16'b0;
    assign data[9435] = ~16'b0;
    assign data[9436] = ~16'b0;
    assign data[9437] = ~16'b0;
    assign data[9438] = ~16'b0;
    assign data[9439] = ~16'b0;
    assign data[9440] = ~16'b0;
    assign data[9441] = ~16'b0;
    assign data[9442] = ~16'b0;
    assign data[9443] = ~16'b0;
    assign data[9444] = ~16'b0;
    assign data[9445] = ~16'b0;
    assign data[9446] = ~16'b0;
    assign data[9447] = ~16'b0;
    assign data[9448] = ~16'b0;
    assign data[9449] = ~16'b0;
    assign data[9450] = ~16'b0;
    assign data[9451] = ~16'b0;
    assign data[9452] = ~16'b0;
    assign data[9453] = ~16'b0;
    assign data[9454] = ~16'b0;
    assign data[9455] = ~16'b0;
    assign data[9456] = ~16'b0;
    assign data[9457] = ~16'b0;
    assign data[9458] = ~16'b0;
    assign data[9459] = ~16'b0;
    assign data[9460] = ~16'b0;
    assign data[9461] = ~16'b0;
    assign data[9462] = ~16'b0;
    assign data[9463] = ~16'b0;
    assign data[9464] = ~16'b0;
    assign data[9465] = ~16'b0;
    assign data[9466] = ~16'b0;
    assign data[9467] = ~16'b0;
    assign data[9468] = ~16'b0;
    assign data[9469] = ~16'b0;
    assign data[9470] = ~16'b0;
    assign data[9471] = ~16'b0;
    assign data[9472] = ~16'b0;
    assign data[9473] = ~16'b0;
    assign data[9474] = ~16'b0;
    assign data[9475] = ~16'b0;
    assign data[9476] = ~16'b0;
    assign data[9477] = ~16'b0;
    assign data[9478] = ~16'b0;
    assign data[9479] = ~16'b0;
    assign data[9480] = ~16'b0;
    assign data[9481] = ~16'b0;
    assign data[9482] = ~16'b0;
    assign data[9483] = ~16'b0;
    assign data[9484] = ~16'b0;
    assign data[9485] = ~16'b0;
    assign data[9486] = ~16'b0;
    assign data[9487] = ~16'b0;
    assign data[9488] = ~16'b0;
    assign data[9489] = ~16'b0;
    assign data[9490] = 16'b0;
    assign data[9491] = 16'b0;
    assign data[9492] = 16'b0;
    assign data[9493] = 16'b0;
    assign data[9494] = 16'b0;
    assign data[9495] = 16'b0;
    assign data[9496] = 16'b0;
    assign data[9497] = 16'b0;
    assign data[9498] = 16'b0;
    assign data[9499] = 16'b0;
    assign data[9500] = 16'b0;
    assign data[9501] = 16'b0;
    assign data[9502] = 16'b0;
    assign data[9503] = 16'b0;
    assign data[9504] = 16'b0;
    assign data[9505] = 16'b0;
    assign data[9506] = 16'b0;
    assign data[9507] = 16'b0;
    assign data[9508] = 16'b0;
    assign data[9509] = 16'b0;
    assign data[9510] = 16'b0;
    assign data[9511] = 16'b0;
    assign data[9512] = ~16'b0;
    assign data[9513] = ~16'b0;
    assign data[9514] = ~16'b0;
    assign data[9515] = ~16'b0;
    assign data[9516] = ~16'b0;
    assign data[9517] = ~16'b0;
    assign data[9518] = ~16'b0;
    assign data[9519] = ~16'b0;
    assign data[9520] = 16'b0;
    assign data[9521] = 16'b0;
    assign data[9522] = ~16'b0;
    assign data[9523] = ~16'b0;
    assign data[9524] = ~16'b0;
    assign data[9525] = ~16'b0;
    assign data[9526] = ~16'b0;
    assign data[9527] = ~16'b0;
    assign data[9528] = ~16'b0;
    assign data[9529] = ~16'b0;
    assign data[9530] = 16'b0;
    assign data[9531] = 16'b0;
    assign data[9532] = ~16'b0;
    assign data[9533] = ~16'b0;
    assign data[9534] = ~16'b0;
    assign data[9535] = ~16'b0;
    assign data[9536] = ~16'b0;
    assign data[9537] = ~16'b0;
    assign data[9538] = ~16'b0;
    assign data[9539] = ~16'b0;
    assign data[9540] = 16'b0;
    assign data[9541] = 16'b0;
    assign data[9542] = ~16'b0;
    assign data[9543] = ~16'b0;
    assign data[9544] = ~16'b0;
    assign data[9545] = ~16'b0;
    assign data[9546] = ~16'b0;
    assign data[9547] = ~16'b0;
    assign data[9548] = ~16'b0;
    assign data[9549] = ~16'b0;
    assign data[9550] = 16'b0;
    assign data[9551] = 16'b0;
    assign data[9552] = ~16'b0;
    assign data[9553] = ~16'b0;
    assign data[9554] = ~16'b0;
    assign data[9555] = ~16'b0;
    assign data[9556] = ~16'b0;
    assign data[9557] = ~16'b0;
    assign data[9558] = ~16'b0;
    assign data[9559] = ~16'b0;
    assign data[9560] = 16'b0;
    assign data[9561] = 16'b0;
    assign data[9562] = ~16'b0;
    assign data[9563] = ~16'b0;
    assign data[9564] = ~16'b0;
    assign data[9565] = ~16'b0;
    assign data[9566] = ~16'b0;
    assign data[9567] = ~16'b0;
    assign data[9568] = ~16'b0;
    assign data[9569] = ~16'b0;
    assign data[9570] = 16'b0;
    assign data[9571] = 16'b0;
    assign data[9572] = ~16'b0;
    assign data[9573] = ~16'b0;
    assign data[9574] = ~16'b0;
    assign data[9575] = ~16'b0;
    assign data[9576] = ~16'b0;
    assign data[9577] = ~16'b0;
    assign data[9578] = ~16'b0;
    assign data[9579] = ~16'b0;
    assign data[9580] = 16'b0;
    assign data[9581] = 16'b0;
    assign data[9582] = ~16'b0;
    assign data[9583] = ~16'b0;
    assign data[9584] = ~16'b0;
    assign data[9585] = ~16'b0;
    assign data[9586] = ~16'b0;
    assign data[9587] = ~16'b0;
    assign data[9588] = ~16'b0;
    assign data[9589] = ~16'b0;
    assign data[9590] = 16'b0;
    assign data[9591] = 16'b0;
    assign data[9592] = ~16'b0;
    assign data[9593] = ~16'b0;
    assign data[9594] = ~16'b0;
    assign data[9595] = ~16'b0;
    assign data[9596] = ~16'b0;
    assign data[9597] = ~16'b0;
    assign data[9598] = ~16'b0;
    assign data[9599] = ~16'b0;
    assign data[9600] = 16'b0;
    assign data[9601] = 16'b0;
    assign data[9602] = ~16'b0;
    assign data[9603] = ~16'b0;
    assign data[9604] = ~16'b0;
    assign data[9605] = ~16'b0;
    assign data[9606] = ~16'b0;
    assign data[9607] = ~16'b0;
    assign data[9608] = ~16'b0;
    assign data[9609] = ~16'b0;
    assign data[9610] = 16'b0;
    assign data[9611] = 16'b0;
    assign data[9612] = ~16'b0;
    assign data[9613] = ~16'b0;
    assign data[9614] = ~16'b0;
    assign data[9615] = ~16'b0;
    assign data[9616] = ~16'b0;
    assign data[9617] = ~16'b0;
    assign data[9618] = ~16'b0;
    assign data[9619] = ~16'b0;
    assign data[9620] = 16'b0;
    assign data[9621] = 16'b0;
    assign data[9622] = ~16'b0;
    assign data[9623] = ~16'b0;
    assign data[9624] = ~16'b0;
    assign data[9625] = ~16'b0;
    assign data[9626] = ~16'b0;
    assign data[9627] = ~16'b0;
    assign data[9628] = ~16'b0;
    assign data[9629] = ~16'b0;
    assign data[9630] = 16'b0;
    assign data[9631] = 16'b0;
    assign data[9632] = ~16'b0;
    assign data[9633] = ~16'b0;
    assign data[9634] = ~16'b0;
    assign data[9635] = ~16'b0;
    assign data[9636] = ~16'b0;
    assign data[9637] = ~16'b0;
    assign data[9638] = ~16'b0;
    assign data[9639] = ~16'b0;
    assign data[9640] = 16'b0;
    assign data[9641] = 16'b0;
    assign data[9642] = ~16'b0;
    assign data[9643] = ~16'b0;
    assign data[9644] = ~16'b0;
    assign data[9645] = ~16'b0;
    assign data[9646] = ~16'b0;
    assign data[9647] = ~16'b0;
    assign data[9648] = ~16'b0;
    assign data[9649] = ~16'b0;
    assign data[9650] = 16'b0;
    assign data[9651] = 16'b0;
    assign data[9652] = ~16'b0;
    assign data[9653] = ~16'b0;
    assign data[9654] = ~16'b0;
    assign data[9655] = ~16'b0;
    assign data[9656] = ~16'b0;
    assign data[9657] = ~16'b0;
    assign data[9658] = ~16'b0;
    assign data[9659] = ~16'b0;
    assign data[9660] = 16'b0;
    assign data[9661] = 16'b0;
    assign data[9662] = ~16'b0;
    assign data[9663] = ~16'b0;
    assign data[9664] = ~16'b0;
    assign data[9665] = ~16'b0;
    assign data[9666] = ~16'b0;
    assign data[9667] = ~16'b0;
    assign data[9668] = ~16'b0;
    assign data[9669] = ~16'b0;
    assign data[9670] = 16'b0;
    assign data[9671] = 16'b0;
    assign data[9672] = ~16'b0;
    assign data[9673] = ~16'b0;
    assign data[9674] = ~16'b0;
    assign data[9675] = ~16'b0;
    assign data[9676] = ~16'b0;
    assign data[9677] = ~16'b0;
    assign data[9678] = ~16'b0;
    assign data[9679] = ~16'b0;
    assign data[9680] = 16'b0;
    assign data[9681] = 16'b0;
    assign data[9682] = ~16'b0;
    assign data[9683] = ~16'b0;
    assign data[9684] = ~16'b0;
    assign data[9685] = ~16'b0;
    assign data[9686] = ~16'b0;
    assign data[9687] = ~16'b0;
    assign data[9688] = ~16'b0;
    assign data[9689] = ~16'b0;
    assign data[9690] = 16'b0;
    assign data[9691] = 16'b0;
    assign data[9692] = ~16'b0;
    assign data[9693] = ~16'b0;
    assign data[9694] = ~16'b0;
    assign data[9695] = ~16'b0;
    assign data[9696] = ~16'b0;
    assign data[9697] = ~16'b0;
    assign data[9698] = ~16'b0;
    assign data[9699] = ~16'b0;
    assign data[9700] = 16'b0;
    assign data[9701] = 16'b0;
    assign data[9702] = ~16'b0;
    assign data[9703] = ~16'b0;
    assign data[9704] = ~16'b0;
    assign data[9705] = ~16'b0;
    assign data[9706] = ~16'b0;
    assign data[9707] = ~16'b0;
    assign data[9708] = ~16'b0;
    assign data[9709] = ~16'b0;
    assign data[9710] = 16'b0;
    assign data[9711] = 16'b0;
    assign data[9712] = ~16'b0;
    assign data[9713] = ~16'b0;
    assign data[9714] = ~16'b0;
    assign data[9715] = ~16'b0;
    assign data[9716] = ~16'b0;
    assign data[9717] = ~16'b0;
    assign data[9718] = ~16'b0;
    assign data[9719] = ~16'b0;
    assign data[9720] = 16'b0;
    assign data[9721] = 16'b0;
    assign data[9722] = ~16'b0;
    assign data[9723] = ~16'b0;
    assign data[9724] = ~16'b0;
    assign data[9725] = ~16'b0;
    assign data[9726] = ~16'b0;
    assign data[9727] = ~16'b0;
    assign data[9728] = ~16'b0;
    assign data[9729] = ~16'b0;
    assign data[9730] = 16'b0;
    assign data[9731] = 16'b0;
    assign data[9732] = ~16'b0;
    assign data[9733] = ~16'b0;
    assign data[9734] = ~16'b0;
    assign data[9735] = ~16'b0;
    assign data[9736] = ~16'b0;
    assign data[9737] = ~16'b0;
    assign data[9738] = ~16'b0;
    assign data[9739] = ~16'b0;
    assign data[9740] = 16'b0;
    assign data[9741] = 16'b0;
    assign data[9742] = ~16'b0;
    assign data[9743] = ~16'b0;
    assign data[9744] = ~16'b0;
    assign data[9745] = ~16'b0;
    assign data[9746] = ~16'b0;
    assign data[9747] = ~16'b0;
    assign data[9748] = ~16'b0;
    assign data[9749] = ~16'b0;
    assign data[9750] = 16'b0;
    assign data[9751] = 16'b0;
    assign data[9752] = ~16'b0;
    assign data[9753] = ~16'b0;
    assign data[9754] = ~16'b0;
    assign data[9755] = ~16'b0;
    assign data[9756] = ~16'b0;
    assign data[9757] = ~16'b0;
    assign data[9758] = ~16'b0;
    assign data[9759] = ~16'b0;
    assign data[9760] = 16'b0;
    assign data[9761] = 16'b0;
    assign data[9762] = ~16'b0;
    assign data[9763] = ~16'b0;
    assign data[9764] = ~16'b0;
    assign data[9765] = ~16'b0;
    assign data[9766] = ~16'b0;
    assign data[9767] = ~16'b0;
    assign data[9768] = ~16'b0;
    assign data[9769] = ~16'b0;
    assign data[9770] = 16'b0;
    assign data[9771] = 16'b0;
    assign data[9772] = ~16'b0;
    assign data[9773] = ~16'b0;
    assign data[9774] = ~16'b0;
    assign data[9775] = ~16'b0;
    assign data[9776] = ~16'b0;
    assign data[9777] = ~16'b0;
    assign data[9778] = ~16'b0;
    assign data[9779] = ~16'b0;
    assign data[9780] = 16'b0;
    assign data[9781] = 16'b0;
    assign data[9782] = ~16'b0;
    assign data[9783] = ~16'b0;
    assign data[9784] = ~16'b0;
    assign data[9785] = ~16'b0;
    assign data[9786] = ~16'b0;
    assign data[9787] = ~16'b0;
    assign data[9788] = ~16'b0;
    assign data[9789] = ~16'b0;
    assign data[9790] = 16'b0;
    assign data[9791] = 16'b0;
    assign data[9792] = ~16'b0;
    assign data[9793] = ~16'b0;
    assign data[9794] = ~16'b0;
    assign data[9795] = ~16'b0;
    assign data[9796] = ~16'b0;
    assign data[9797] = ~16'b0;
    assign data[9798] = ~16'b0;
    assign data[9799] = ~16'b0;
    assign data[9800] = 16'b0;
    assign data[9801] = 16'b0;
    assign data[9802] = ~16'b0;
    assign data[9803] = ~16'b0;
    assign data[9804] = ~16'b0;
    assign data[9805] = ~16'b0;
    assign data[9806] = ~16'b0;
    assign data[9807] = ~16'b0;
    assign data[9808] = ~16'b0;
    assign data[9809] = ~16'b0;
    assign data[9810] = 16'b0;
    assign data[9811] = 16'b0;
    assign data[9812] = ~16'b0;
    assign data[9813] = ~16'b0;
    assign data[9814] = ~16'b0;
    assign data[9815] = ~16'b0;
    assign data[9816] = ~16'b0;
    assign data[9817] = ~16'b0;
    assign data[9818] = ~16'b0;
    assign data[9819] = ~16'b0;
    assign data[9820] = 16'b0;
    assign data[9821] = 16'b0;
    assign data[9822] = ~16'b0;
    assign data[9823] = ~16'b0;
    assign data[9824] = ~16'b0;
    assign data[9825] = ~16'b0;
    assign data[9826] = ~16'b0;
    assign data[9827] = ~16'b0;
    assign data[9828] = ~16'b0;
    assign data[9829] = ~16'b0;
    assign data[9830] = 16'b0;
    assign data[9831] = 16'b0;
    assign data[9832] = ~16'b0;
    assign data[9833] = ~16'b0;
    assign data[9834] = ~16'b0;
    assign data[9835] = ~16'b0;
    assign data[9836] = ~16'b0;
    assign data[9837] = ~16'b0;
    assign data[9838] = ~16'b0;
    assign data[9839] = ~16'b0;
    assign data[9840] = 16'b0;
    assign data[9841] = 16'b0;
    assign data[9842] = 16'b0;
    assign data[9843] = 16'b0;
    assign data[9844] = 16'b0;
    assign data[9845] = 16'b0;
    assign data[9846] = 16'b0;
    assign data[9847] = 16'b0;
    assign data[9848] = 16'b0;
    assign data[9849] = 16'b0;
    assign data[9850] = 16'b0;
    assign data[9851] = 16'b0;
    assign data[9852] = 16'b0;
    assign data[9853] = 16'b0;
    assign data[9854] = 16'b0;
    assign data[9855] = 16'b0;
    assign data[9856] = 16'b0;
    assign data[9857] = 16'b0;
    assign data[9858] = 16'b0;
    assign data[9859] = 16'b0;
    assign data[9860] = ~16'b0;
    assign data[9861] = ~16'b0;
    assign data[9862] = ~16'b0;
    assign data[9863] = ~16'b0;
    assign data[9864] = ~16'b0;
    assign data[9865] = ~16'b0;
    assign data[9866] = ~16'b0;
    assign data[9867] = ~16'b0;
    assign data[9868] = ~16'b0;
    assign data[9869] = ~16'b0;
    assign data[9870] = ~16'b0;
    assign data[9871] = ~16'b0;
    assign data[9872] = ~16'b0;
    assign data[9873] = ~16'b0;
    assign data[9874] = ~16'b0;
    assign data[9875] = ~16'b0;
    assign data[9876] = ~16'b0;
    assign data[9877] = ~16'b0;
    assign data[9878] = ~16'b0;
    assign data[9879] = ~16'b0;
    assign data[9880] = ~16'b0;
    assign data[9881] = ~16'b0;
    assign data[9882] = ~16'b0;
    assign data[9883] = ~16'b0;
    assign data[9884] = ~16'b0;
    assign data[9885] = ~16'b0;
    assign data[9886] = ~16'b0;
    assign data[9887] = ~16'b0;
    assign data[9888] = ~16'b0;
    assign data[9889] = ~16'b0;
    assign data[9890] = ~16'b0;
    assign data[9891] = ~16'b0;
    assign data[9892] = ~16'b0;
    assign data[9893] = ~16'b0;
    assign data[9894] = ~16'b0;
    assign data[9895] = ~16'b0;
    assign data[9896] = ~16'b0;
    assign data[9897] = ~16'b0;
    assign data[9898] = ~16'b0;
    assign data[9899] = ~16'b0;
    assign data[9900] = ~16'b0;
    assign data[9901] = ~16'b0;
    assign data[9902] = ~16'b0;
    assign data[9903] = ~16'b0;
    assign data[9904] = ~16'b0;
    assign data[9905] = ~16'b0;
    assign data[9906] = ~16'b0;
    assign data[9907] = ~16'b0;
    assign data[9908] = ~16'b0;
    assign data[9909] = ~16'b0;
    assign data[9910] = ~16'b0;
    assign data[9911] = ~16'b0;
    assign data[9912] = ~16'b0;
    assign data[9913] = ~16'b0;
    assign data[9914] = ~16'b0;
    assign data[9915] = ~16'b0;
    assign data[9916] = ~16'b0;
    assign data[9917] = ~16'b0;
    assign data[9918] = ~16'b0;
    assign data[9919] = ~16'b0;
    assign data[9920] = ~16'b0;
    assign data[9921] = ~16'b0;
    assign data[9922] = ~16'b0;
    assign data[9923] = ~16'b0;
    assign data[9924] = ~16'b0;
    assign data[9925] = ~16'b0;
    assign data[9926] = ~16'b0;
    assign data[9927] = ~16'b0;
    assign data[9928] = ~16'b0;
    assign data[9929] = ~16'b0;
    assign data[9930] = ~16'b0;
    assign data[9931] = ~16'b0;
    assign data[9932] = ~16'b0;
    assign data[9933] = ~16'b0;
    assign data[9934] = ~16'b0;
    assign data[9935] = ~16'b0;
    assign data[9936] = ~16'b0;
    assign data[9937] = ~16'b0;
    assign data[9938] = ~16'b0;
    assign data[9939] = ~16'b0;
    assign data[9940] = ~16'b0;
    assign data[9941] = ~16'b0;
    assign data[9942] = ~16'b0;
    assign data[9943] = ~16'b0;
    assign data[9944] = ~16'b0;
    assign data[9945] = ~16'b0;
    assign data[9946] = ~16'b0;
    assign data[9947] = ~16'b0;
    assign data[9948] = ~16'b0;
    assign data[9949] = ~16'b0;
    assign data[9950] = ~16'b0;
    assign data[9951] = ~16'b0;
    assign data[9952] = ~16'b0;
    assign data[9953] = ~16'b0;
    assign data[9954] = ~16'b0;
    assign data[9955] = ~16'b0;
    assign data[9956] = ~16'b0;
    assign data[9957] = ~16'b0;
    assign data[9958] = ~16'b0;
    assign data[9959] = ~16'b0;
    assign data[9960] = ~16'b0;
    assign data[9961] = ~16'b0;
    assign data[9962] = ~16'b0;
    assign data[9963] = ~16'b0;
    assign data[9964] = ~16'b0;
    assign data[9965] = ~16'b0;
    assign data[9966] = ~16'b0;
    assign data[9967] = ~16'b0;
    assign data[9968] = ~16'b0;
    assign data[9969] = ~16'b0;
    assign data[9970] = ~16'b0;
    assign data[9971] = ~16'b0;
    assign data[9972] = ~16'b0;
    assign data[9973] = ~16'b0;
    assign data[9974] = ~16'b0;
    assign data[9975] = ~16'b0;
    assign data[9976] = ~16'b0;
    assign data[9977] = ~16'b0;
    assign data[9978] = ~16'b0;
    assign data[9979] = ~16'b0;
    assign data[9980] = ~16'b0;
    assign data[9981] = ~16'b0;
    assign data[9982] = ~16'b0;
    assign data[9983] = ~16'b0;
    assign data[9984] = ~16'b0;
    assign data[9985] = ~16'b0;
    assign data[9986] = ~16'b0;
    assign data[9987] = ~16'b0;
    assign data[9988] = ~16'b0;
    assign data[9989] = ~16'b0;
    assign data[9990] = ~16'b0;
    assign data[9991] = ~16'b0;
    assign data[9992] = ~16'b0;
    assign data[9993] = ~16'b0;
    assign data[9994] = ~16'b0;
    assign data[9995] = ~16'b0;
    assign data[9996] = ~16'b0;
    assign data[9997] = ~16'b0;
    assign data[9998] = ~16'b0;
    assign data[9999] = ~16'b0;
    assign data[10000] = ~16'b0;
    assign data[10001] = ~16'b0;
    assign data[10002] = ~16'b0;
    assign data[10003] = ~16'b0;
    assign data[10004] = ~16'b0;
    assign data[10005] = ~16'b0;
    assign data[10006] = ~16'b0;
    assign data[10007] = ~16'b0;
    assign data[10008] = ~16'b0;
    assign data[10009] = ~16'b0;
    assign data[10010] = ~16'b0;
    assign data[10011] = ~16'b0;
    assign data[10012] = ~16'b0;
    assign data[10013] = ~16'b0;
    assign data[10014] = ~16'b0;
    assign data[10015] = ~16'b0;
    assign data[10016] = ~16'b0;
    assign data[10017] = ~16'b0;
    assign data[10018] = ~16'b0;
    assign data[10019] = ~16'b0;
    assign data[10020] = ~16'b0;
    assign data[10021] = ~16'b0;
    assign data[10022] = ~16'b0;
    assign data[10023] = ~16'b0;
    assign data[10024] = ~16'b0;
    assign data[10025] = ~16'b0;
    assign data[10026] = ~16'b0;
    assign data[10027] = ~16'b0;
    assign data[10028] = ~16'b0;
    assign data[10029] = ~16'b0;
    assign data[10030] = ~16'b0;
    assign data[10031] = ~16'b0;
    assign data[10032] = ~16'b0;
    assign data[10033] = ~16'b0;
    assign data[10034] = ~16'b0;
    assign data[10035] = ~16'b0;
    assign data[10036] = ~16'b0;
    assign data[10037] = ~16'b0;
    assign data[10038] = ~16'b0;
    assign data[10039] = ~16'b0;
    assign data[10040] = ~16'b0;
    assign data[10041] = ~16'b0;
    assign data[10042] = ~16'b0;
    assign data[10043] = ~16'b0;
    assign data[10044] = ~16'b0;
    assign data[10045] = ~16'b0;
    assign data[10046] = ~16'b0;
    assign data[10047] = ~16'b0;
    assign data[10048] = ~16'b0;
    assign data[10049] = ~16'b0;
    assign data[10050] = ~16'b0;
    assign data[10051] = ~16'b0;
    assign data[10052] = ~16'b0;
    assign data[10053] = ~16'b0;
    assign data[10054] = ~16'b0;
    assign data[10055] = ~16'b0;
    assign data[10056] = ~16'b0;
    assign data[10057] = ~16'b0;
    assign data[10058] = ~16'b0;
    assign data[10059] = ~16'b0;
    assign data[10060] = ~16'b0;
    assign data[10061] = ~16'b0;
    assign data[10062] = ~16'b0;
    assign data[10063] = ~16'b0;
    assign data[10064] = ~16'b0;
    assign data[10065] = ~16'b0;
    assign data[10066] = ~16'b0;
    assign data[10067] = ~16'b0;
    assign data[10068] = ~16'b0;
    assign data[10069] = ~16'b0;
    assign data[10070] = 16'b0;
    assign data[10071] = 16'b0;
    assign data[10072] = 16'b0;
    assign data[10073] = 16'b0;
    assign data[10074] = 16'b0;
    assign data[10075] = 16'b0;
    assign data[10076] = 16'b0;
    assign data[10077] = 16'b0;
    assign data[10078] = 16'b0;
    assign data[10079] = 16'b0;
    assign data[10080] = 16'b0;
    assign data[10081] = 16'b0;
    assign data[10082] = 16'b0;
    assign data[10083] = 16'b0;
    assign data[10084] = 16'b0;
    assign data[10085] = 16'b0;
    assign data[10086] = 16'b0;
    assign data[10087] = 16'b0;
    assign data[10088] = 16'b0;
    assign data[10089] = 16'b0;
    assign data[10090] = 16'b0;
    assign data[10091] = 16'b0;
    assign data[10092] = ~16'b0;
    assign data[10093] = ~16'b0;
    assign data[10094] = ~16'b0;
    assign data[10095] = ~16'b0;
    assign data[10096] = ~16'b0;
    assign data[10097] = ~16'b0;
    assign data[10098] = ~16'b0;
    assign data[10099] = ~16'b0;
    assign data[10100] = 16'b0;
    assign data[10101] = 16'b0;
    assign data[10102] = ~16'b0;
    assign data[10103] = ~16'b0;
    assign data[10104] = ~16'b0;
    assign data[10105] = ~16'b0;
    assign data[10106] = ~16'b0;
    assign data[10107] = ~16'b0;
    assign data[10108] = ~16'b0;
    assign data[10109] = ~16'b0;
    assign data[10110] = 16'b0;
    assign data[10111] = 16'b0;
    assign data[10112] = ~16'b0;
    assign data[10113] = ~16'b0;
    assign data[10114] = ~16'b0;
    assign data[10115] = ~16'b0;
    assign data[10116] = ~16'b0;
    assign data[10117] = ~16'b0;
    assign data[10118] = ~16'b0;
    assign data[10119] = ~16'b0;
    assign data[10120] = 16'b0;
    assign data[10121] = 16'b0;
    assign data[10122] = ~16'b0;
    assign data[10123] = ~16'b0;
    assign data[10124] = ~16'b0;
    assign data[10125] = ~16'b0;
    assign data[10126] = ~16'b0;
    assign data[10127] = ~16'b0;
    assign data[10128] = ~16'b0;
    assign data[10129] = ~16'b0;
    assign data[10130] = 16'b0;
    assign data[10131] = 16'b0;
    assign data[10132] = ~16'b0;
    assign data[10133] = ~16'b0;
    assign data[10134] = ~16'b0;
    assign data[10135] = ~16'b0;
    assign data[10136] = ~16'b0;
    assign data[10137] = ~16'b0;
    assign data[10138] = ~16'b0;
    assign data[10139] = ~16'b0;
    assign data[10140] = 16'b0;
    assign data[10141] = 16'b0;
    assign data[10142] = ~16'b0;
    assign data[10143] = ~16'b0;
    assign data[10144] = ~16'b0;
    assign data[10145] = ~16'b0;
    assign data[10146] = ~16'b0;
    assign data[10147] = ~16'b0;
    assign data[10148] = ~16'b0;
    assign data[10149] = ~16'b0;
    assign data[10150] = 16'b0;
    assign data[10151] = 16'b0;
    assign data[10152] = ~16'b0;
    assign data[10153] = ~16'b0;
    assign data[10154] = ~16'b0;
    assign data[10155] = ~16'b0;
    assign data[10156] = ~16'b0;
    assign data[10157] = ~16'b0;
    assign data[10158] = ~16'b0;
    assign data[10159] = ~16'b0;
    assign data[10160] = 16'b0;
    assign data[10161] = 16'b0;
    assign data[10162] = ~16'b0;
    assign data[10163] = ~16'b0;
    assign data[10164] = ~16'b0;
    assign data[10165] = ~16'b0;
    assign data[10166] = ~16'b0;
    assign data[10167] = ~16'b0;
    assign data[10168] = ~16'b0;
    assign data[10169] = ~16'b0;
    assign data[10170] = 16'b0;
    assign data[10171] = 16'b0;
    assign data[10172] = ~16'b0;
    assign data[10173] = ~16'b0;
    assign data[10174] = ~16'b0;
    assign data[10175] = ~16'b0;
    assign data[10176] = ~16'b0;
    assign data[10177] = ~16'b0;
    assign data[10178] = ~16'b0;
    assign data[10179] = ~16'b0;
    assign data[10180] = 16'b0;
    assign data[10181] = 16'b0;
    assign data[10182] = ~16'b0;
    assign data[10183] = ~16'b0;
    assign data[10184] = ~16'b0;
    assign data[10185] = ~16'b0;
    assign data[10186] = ~16'b0;
    assign data[10187] = ~16'b0;
    assign data[10188] = ~16'b0;
    assign data[10189] = ~16'b0;
    assign data[10190] = 16'b0;
    assign data[10191] = 16'b0;
    assign data[10192] = ~16'b0;
    assign data[10193] = ~16'b0;
    assign data[10194] = ~16'b0;
    assign data[10195] = ~16'b0;
    assign data[10196] = ~16'b0;
    assign data[10197] = ~16'b0;
    assign data[10198] = ~16'b0;
    assign data[10199] = ~16'b0;
    assign data[10200] = 16'b0;
    assign data[10201] = 16'b0;
    assign data[10202] = ~16'b0;
    assign data[10203] = ~16'b0;
    assign data[10204] = ~16'b0;
    assign data[10205] = ~16'b0;
    assign data[10206] = ~16'b0;
    assign data[10207] = ~16'b0;
    assign data[10208] = ~16'b0;
    assign data[10209] = ~16'b0;
    assign data[10210] = 16'b0;
    assign data[10211] = 16'b0;
    assign data[10212] = ~16'b0;
    assign data[10213] = ~16'b0;
    assign data[10214] = ~16'b0;
    assign data[10215] = ~16'b0;
    assign data[10216] = ~16'b0;
    assign data[10217] = ~16'b0;
    assign data[10218] = ~16'b0;
    assign data[10219] = ~16'b0;
    assign data[10220] = 16'b0;
    assign data[10221] = 16'b0;
    assign data[10222] = ~16'b0;
    assign data[10223] = ~16'b0;
    assign data[10224] = ~16'b0;
    assign data[10225] = ~16'b0;
    assign data[10226] = ~16'b0;
    assign data[10227] = ~16'b0;
    assign data[10228] = ~16'b0;
    assign data[10229] = ~16'b0;
    assign data[10230] = 16'b0;
    assign data[10231] = 16'b0;
    assign data[10232] = ~16'b0;
    assign data[10233] = ~16'b0;
    assign data[10234] = ~16'b0;
    assign data[10235] = ~16'b0;
    assign data[10236] = ~16'b0;
    assign data[10237] = ~16'b0;
    assign data[10238] = ~16'b0;
    assign data[10239] = ~16'b0;
    assign data[10240] = 16'b0;
    assign data[10241] = 16'b0;
    assign data[10242] = ~16'b0;
    assign data[10243] = ~16'b0;
    assign data[10244] = ~16'b0;
    assign data[10245] = ~16'b0;
    assign data[10246] = ~16'b0;
    assign data[10247] = ~16'b0;
    assign data[10248] = ~16'b0;
    assign data[10249] = ~16'b0;
    assign data[10250] = 16'b0;
    assign data[10251] = 16'b0;
    assign data[10252] = ~16'b0;
    assign data[10253] = ~16'b0;
    assign data[10254] = ~16'b0;
    assign data[10255] = ~16'b0;
    assign data[10256] = ~16'b0;
    assign data[10257] = ~16'b0;
    assign data[10258] = ~16'b0;
    assign data[10259] = ~16'b0;
    assign data[10260] = 16'b0;
    assign data[10261] = 16'b0;
    assign data[10262] = ~16'b0;
    assign data[10263] = ~16'b0;
    assign data[10264] = ~16'b0;
    assign data[10265] = ~16'b0;
    assign data[10266] = ~16'b0;
    assign data[10267] = ~16'b0;
    assign data[10268] = ~16'b0;
    assign data[10269] = ~16'b0;
    assign data[10270] = 16'b0;
    assign data[10271] = 16'b0;
    assign data[10272] = ~16'b0;
    assign data[10273] = ~16'b0;
    assign data[10274] = ~16'b0;
    assign data[10275] = ~16'b0;
    assign data[10276] = ~16'b0;
    assign data[10277] = ~16'b0;
    assign data[10278] = ~16'b0;
    assign data[10279] = ~16'b0;
    assign data[10280] = 16'b0;
    assign data[10281] = 16'b0;
    assign data[10282] = ~16'b0;
    assign data[10283] = ~16'b0;
    assign data[10284] = ~16'b0;
    assign data[10285] = ~16'b0;
    assign data[10286] = ~16'b0;
    assign data[10287] = ~16'b0;
    assign data[10288] = ~16'b0;
    assign data[10289] = ~16'b0;
    assign data[10290] = 16'b0;
    assign data[10291] = 16'b0;
    assign data[10292] = ~16'b0;
    assign data[10293] = ~16'b0;
    assign data[10294] = ~16'b0;
    assign data[10295] = ~16'b0;
    assign data[10296] = ~16'b0;
    assign data[10297] = ~16'b0;
    assign data[10298] = ~16'b0;
    assign data[10299] = ~16'b0;
    assign data[10300] = 16'b0;
    assign data[10301] = 16'b0;
    assign data[10302] = ~16'b0;
    assign data[10303] = ~16'b0;
    assign data[10304] = ~16'b0;
    assign data[10305] = ~16'b0;
    assign data[10306] = ~16'b0;
    assign data[10307] = ~16'b0;
    assign data[10308] = ~16'b0;
    assign data[10309] = ~16'b0;
    assign data[10310] = 16'b0;
    assign data[10311] = 16'b0;
    assign data[10312] = ~16'b0;
    assign data[10313] = ~16'b0;
    assign data[10314] = ~16'b0;
    assign data[10315] = ~16'b0;
    assign data[10316] = ~16'b0;
    assign data[10317] = ~16'b0;
    assign data[10318] = ~16'b0;
    assign data[10319] = ~16'b0;
    assign data[10320] = 16'b0;
    assign data[10321] = 16'b0;
    assign data[10322] = ~16'b0;
    assign data[10323] = ~16'b0;
    assign data[10324] = ~16'b0;
    assign data[10325] = ~16'b0;
    assign data[10326] = ~16'b0;
    assign data[10327] = ~16'b0;
    assign data[10328] = ~16'b0;
    assign data[10329] = ~16'b0;
    assign data[10330] = 16'b0;
    assign data[10331] = 16'b0;
    assign data[10332] = ~16'b0;
    assign data[10333] = ~16'b0;
    assign data[10334] = ~16'b0;
    assign data[10335] = ~16'b0;
    assign data[10336] = ~16'b0;
    assign data[10337] = ~16'b0;
    assign data[10338] = ~16'b0;
    assign data[10339] = ~16'b0;
    assign data[10340] = 16'b0;
    assign data[10341] = 16'b0;
    assign data[10342] = ~16'b0;
    assign data[10343] = ~16'b0;
    assign data[10344] = ~16'b0;
    assign data[10345] = ~16'b0;
    assign data[10346] = ~16'b0;
    assign data[10347] = ~16'b0;
    assign data[10348] = ~16'b0;
    assign data[10349] = ~16'b0;
    assign data[10350] = 16'b0;
    assign data[10351] = 16'b0;
    assign data[10352] = 16'b0;
    assign data[10353] = 16'b0;
    assign data[10354] = 16'b0;
    assign data[10355] = 16'b0;
    assign data[10356] = 16'b0;
    assign data[10357] = 16'b0;
    assign data[10358] = 16'b0;
    assign data[10359] = 16'b0;
    assign data[10360] = 16'b0;
    assign data[10361] = 16'b0;
    assign data[10362] = 16'b0;
    assign data[10363] = 16'b0;
    assign data[10364] = 16'b0;
    assign data[10365] = 16'b0;
    assign data[10366] = 16'b0;
    assign data[10367] = 16'b0;
    assign data[10368] = 16'b0;
    assign data[10369] = 16'b0;
    assign data[10370] = ~16'b0;
    assign data[10371] = ~16'b0;
    assign data[10372] = ~16'b0;
    assign data[10373] = ~16'b0;
    assign data[10374] = ~16'b0;
    assign data[10375] = ~16'b0;
    assign data[10376] = ~16'b0;
    assign data[10377] = ~16'b0;
    assign data[10378] = ~16'b0;
    assign data[10379] = ~16'b0;
    assign data[10380] = ~16'b0;
    assign data[10381] = ~16'b0;
    assign data[10382] = ~16'b0;
    assign data[10383] = ~16'b0;
    assign data[10384] = ~16'b0;
    assign data[10385] = ~16'b0;
    assign data[10386] = ~16'b0;
    assign data[10387] = ~16'b0;
    assign data[10388] = ~16'b0;
    assign data[10389] = ~16'b0;
    assign data[10390] = ~16'b0;
    assign data[10391] = ~16'b0;
    assign data[10392] = ~16'b0;
    assign data[10393] = ~16'b0;
    assign data[10394] = ~16'b0;
    assign data[10395] = ~16'b0;
    assign data[10396] = ~16'b0;
    assign data[10397] = ~16'b0;
    assign data[10398] = ~16'b0;
    assign data[10399] = ~16'b0;
    assign data[10400] = ~16'b0;
    assign data[10401] = ~16'b0;
    assign data[10402] = ~16'b0;
    assign data[10403] = ~16'b0;
    assign data[10404] = ~16'b0;
    assign data[10405] = ~16'b0;
    assign data[10406] = ~16'b0;
    assign data[10407] = ~16'b0;
    assign data[10408] = ~16'b0;
    assign data[10409] = ~16'b0;
    assign data[10410] = ~16'b0;
    assign data[10411] = ~16'b0;
    assign data[10412] = ~16'b0;
    assign data[10413] = ~16'b0;
    assign data[10414] = ~16'b0;
    assign data[10415] = ~16'b0;
    assign data[10416] = ~16'b0;
    assign data[10417] = ~16'b0;
    assign data[10418] = ~16'b0;
    assign data[10419] = ~16'b0;
    assign data[10420] = ~16'b0;
    assign data[10421] = ~16'b0;
    assign data[10422] = ~16'b0;
    assign data[10423] = ~16'b0;
    assign data[10424] = ~16'b0;
    assign data[10425] = ~16'b0;
    assign data[10426] = ~16'b0;
    assign data[10427] = ~16'b0;
    assign data[10428] = ~16'b0;
    assign data[10429] = ~16'b0;
    assign data[10430] = ~16'b0;
    assign data[10431] = ~16'b0;
    assign data[10432] = ~16'b0;
    assign data[10433] = ~16'b0;
    assign data[10434] = ~16'b0;
    assign data[10435] = ~16'b0;
    assign data[10436] = ~16'b0;
    assign data[10437] = ~16'b0;
    assign data[10438] = ~16'b0;
    assign data[10439] = ~16'b0;
    assign data[10440] = ~16'b0;
    assign data[10441] = ~16'b0;
    assign data[10442] = ~16'b0;
    assign data[10443] = ~16'b0;
    assign data[10444] = ~16'b0;
    assign data[10445] = ~16'b0;
    assign data[10446] = ~16'b0;
    assign data[10447] = ~16'b0;
    assign data[10448] = ~16'b0;
    assign data[10449] = ~16'b0;
    assign data[10450] = ~16'b0;
    assign data[10451] = ~16'b0;
    assign data[10452] = ~16'b0;
    assign data[10453] = ~16'b0;
    assign data[10454] = ~16'b0;
    assign data[10455] = ~16'b0;
    assign data[10456] = ~16'b0;
    assign data[10457] = ~16'b0;
    assign data[10458] = ~16'b0;
    assign data[10459] = ~16'b0;
    assign data[10460] = ~16'b0;
    assign data[10461] = ~16'b0;
    assign data[10462] = ~16'b0;
    assign data[10463] = ~16'b0;
    assign data[10464] = ~16'b0;
    assign data[10465] = ~16'b0;
    assign data[10466] = ~16'b0;
    assign data[10467] = ~16'b0;
    assign data[10468] = ~16'b0;
    assign data[10469] = ~16'b0;
    assign data[10470] = ~16'b0;
    assign data[10471] = ~16'b0;
    assign data[10472] = ~16'b0;
    assign data[10473] = ~16'b0;
    assign data[10474] = ~16'b0;
    assign data[10475] = ~16'b0;
    assign data[10476] = ~16'b0;
    assign data[10477] = ~16'b0;
    assign data[10478] = ~16'b0;
    assign data[10479] = ~16'b0;
    assign data[10480] = ~16'b0;
    assign data[10481] = ~16'b0;
    assign data[10482] = ~16'b0;
    assign data[10483] = ~16'b0;
    assign data[10484] = ~16'b0;
    assign data[10485] = ~16'b0;
    assign data[10486] = ~16'b0;
    assign data[10487] = ~16'b0;
    assign data[10488] = ~16'b0;
    assign data[10489] = ~16'b0;
    assign data[10490] = ~16'b0;
    assign data[10491] = ~16'b0;
    assign data[10492] = ~16'b0;
    assign data[10493] = ~16'b0;
    assign data[10494] = ~16'b0;
    assign data[10495] = ~16'b0;
    assign data[10496] = ~16'b0;
    assign data[10497] = ~16'b0;
    assign data[10498] = ~16'b0;
    assign data[10499] = ~16'b0;
    assign data[10500] = ~16'b0;
    assign data[10501] = ~16'b0;
    assign data[10502] = ~16'b0;
    assign data[10503] = ~16'b0;
    assign data[10504] = ~16'b0;
    assign data[10505] = ~16'b0;
    assign data[10506] = ~16'b0;
    assign data[10507] = ~16'b0;
    assign data[10508] = ~16'b0;
    assign data[10509] = ~16'b0;
    assign data[10510] = ~16'b0;
    assign data[10511] = ~16'b0;
    assign data[10512] = ~16'b0;
    assign data[10513] = ~16'b0;
    assign data[10514] = ~16'b0;
    assign data[10515] = ~16'b0;
    assign data[10516] = ~16'b0;
    assign data[10517] = ~16'b0;
    assign data[10518] = ~16'b0;
    assign data[10519] = ~16'b0;
    assign data[10520] = ~16'b0;
    assign data[10521] = ~16'b0;
    assign data[10522] = ~16'b0;
    assign data[10523] = ~16'b0;
    assign data[10524] = ~16'b0;
    assign data[10525] = ~16'b0;
    assign data[10526] = ~16'b0;
    assign data[10527] = ~16'b0;
    assign data[10528] = ~16'b0;
    assign data[10529] = ~16'b0;
    assign data[10530] = ~16'b0;
    assign data[10531] = ~16'b0;
    assign data[10532] = ~16'b0;
    assign data[10533] = ~16'b0;
    assign data[10534] = ~16'b0;
    assign data[10535] = ~16'b0;
    assign data[10536] = ~16'b0;
    assign data[10537] = ~16'b0;
    assign data[10538] = ~16'b0;
    assign data[10539] = ~16'b0;
    assign data[10540] = ~16'b0;
    assign data[10541] = ~16'b0;
    assign data[10542] = ~16'b0;
    assign data[10543] = ~16'b0;
    assign data[10544] = ~16'b0;
    assign data[10545] = ~16'b0;
    assign data[10546] = ~16'b0;
    assign data[10547] = ~16'b0;
    assign data[10548] = ~16'b0;
    assign data[10549] = ~16'b0;
    assign data[10550] = ~16'b0;
    assign data[10551] = ~16'b0;
    assign data[10552] = ~16'b0;
    assign data[10553] = ~16'b0;
    assign data[10554] = ~16'b0;
    assign data[10555] = ~16'b0;
    assign data[10556] = ~16'b0;
    assign data[10557] = ~16'b0;
    assign data[10558] = ~16'b0;
    assign data[10559] = ~16'b0;
    assign data[10560] = ~16'b0;
    assign data[10561] = ~16'b0;
    assign data[10562] = ~16'b0;
    assign data[10563] = ~16'b0;
    assign data[10564] = ~16'b0;
    assign data[10565] = ~16'b0;
    assign data[10566] = ~16'b0;
    assign data[10567] = ~16'b0;
    assign data[10568] = ~16'b0;
    assign data[10569] = ~16'b0;
    assign data[10570] = ~16'b0;
    assign data[10571] = ~16'b0;
    assign data[10572] = ~16'b0;
    assign data[10573] = ~16'b0;
    assign data[10574] = ~16'b0;
    assign data[10575] = ~16'b0;
    assign data[10576] = ~16'b0;
    assign data[10577] = ~16'b0;
    assign data[10578] = ~16'b0;
    assign data[10579] = ~16'b0;
    assign data[10580] = ~16'b0;
    assign data[10581] = ~16'b0;
    assign data[10582] = ~16'b0;
    assign data[10583] = ~16'b0;
    assign data[10584] = ~16'b0;
    assign data[10585] = ~16'b0;
    assign data[10586] = ~16'b0;
    assign data[10587] = ~16'b0;
    assign data[10588] = ~16'b0;
    assign data[10589] = ~16'b0;
    assign data[10590] = ~16'b0;
    assign data[10591] = ~16'b0;
    assign data[10592] = ~16'b0;
    assign data[10593] = ~16'b0;
    assign data[10594] = ~16'b0;
    assign data[10595] = ~16'b0;
    assign data[10596] = ~16'b0;
    assign data[10597] = ~16'b0;
    assign data[10598] = ~16'b0;
    assign data[10599] = ~16'b0;
    assign data[10600] = ~16'b0;
    assign data[10601] = ~16'b0;
    assign data[10602] = ~16'b0;
    assign data[10603] = ~16'b0;
    assign data[10604] = ~16'b0;
    assign data[10605] = ~16'b0;
    assign data[10606] = ~16'b0;
    assign data[10607] = ~16'b0;
    assign data[10608] = ~16'b0;
    assign data[10609] = ~16'b0;
    assign data[10610] = 16'b0;
    assign data[10611] = 16'b0;
    assign data[10612] = 16'b0;
    assign data[10613] = 16'b0;
    assign data[10614] = 16'b0;
    assign data[10615] = 16'b0;
    assign data[10616] = 16'b0;
    assign data[10617] = 16'b0;
    assign data[10618] = 16'b0;
    assign data[10619] = 16'b0;
    assign data[10620] = 16'b0;
    assign data[10621] = 16'b0;
    assign data[10622] = 16'b0;
    assign data[10623] = 16'b0;
    assign data[10624] = 16'b0;
    assign data[10625] = 16'b0;
    assign data[10626] = 16'b0;
    assign data[10627] = 16'b0;
    assign data[10628] = 16'b0;
    assign data[10629] = 16'b0;
    assign data[10630] = 16'b0;
    assign data[10631] = 16'b0;
    assign data[10632] = ~16'b0;
    assign data[10633] = ~16'b0;
    assign data[10634] = ~16'b0;
    assign data[10635] = ~16'b0;
    assign data[10636] = ~16'b0;
    assign data[10637] = ~16'b0;
    assign data[10638] = ~16'b0;
    assign data[10639] = ~16'b0;
    assign data[10640] = 16'b0;
    assign data[10641] = 16'b0;
    assign data[10642] = ~16'b0;
    assign data[10643] = ~16'b0;
    assign data[10644] = ~16'b0;
    assign data[10645] = ~16'b0;
    assign data[10646] = ~16'b0;
    assign data[10647] = ~16'b0;
    assign data[10648] = ~16'b0;
    assign data[10649] = ~16'b0;
    assign data[10650] = 16'b0;
    assign data[10651] = 16'b0;
    assign data[10652] = ~16'b0;
    assign data[10653] = ~16'b0;
    assign data[10654] = ~16'b0;
    assign data[10655] = ~16'b0;
    assign data[10656] = ~16'b0;
    assign data[10657] = ~16'b0;
    assign data[10658] = ~16'b0;
    assign data[10659] = ~16'b0;
    assign data[10660] = 16'b0;
    assign data[10661] = 16'b0;
    assign data[10662] = ~16'b0;
    assign data[10663] = ~16'b0;
    assign data[10664] = ~16'b0;
    assign data[10665] = ~16'b0;
    assign data[10666] = ~16'b0;
    assign data[10667] = ~16'b0;
    assign data[10668] = ~16'b0;
    assign data[10669] = ~16'b0;
    assign data[10670] = 16'b0;
    assign data[10671] = 16'b0;
    assign data[10672] = ~16'b0;
    assign data[10673] = ~16'b0;
    assign data[10674] = ~16'b0;
    assign data[10675] = ~16'b0;
    assign data[10676] = ~16'b0;
    assign data[10677] = ~16'b0;
    assign data[10678] = ~16'b0;
    assign data[10679] = ~16'b0;
    assign data[10680] = 16'b0;
    assign data[10681] = 16'b0;
    assign data[10682] = ~16'b0;
    assign data[10683] = ~16'b0;
    assign data[10684] = ~16'b0;
    assign data[10685] = ~16'b0;
    assign data[10686] = ~16'b0;
    assign data[10687] = ~16'b0;
    assign data[10688] = ~16'b0;
    assign data[10689] = ~16'b0;
    assign data[10690] = 16'b0;
    assign data[10691] = 16'b0;
    assign data[10692] = ~16'b0;
    assign data[10693] = ~16'b0;
    assign data[10694] = ~16'b0;
    assign data[10695] = ~16'b0;
    assign data[10696] = ~16'b0;
    assign data[10697] = ~16'b0;
    assign data[10698] = ~16'b0;
    assign data[10699] = ~16'b0;
    assign data[10700] = 16'b0;
    assign data[10701] = 16'b0;
    assign data[10702] = ~16'b0;
    assign data[10703] = ~16'b0;
    assign data[10704] = ~16'b0;
    assign data[10705] = ~16'b0;
    assign data[10706] = ~16'b0;
    assign data[10707] = ~16'b0;
    assign data[10708] = ~16'b0;
    assign data[10709] = ~16'b0;
    assign data[10710] = 16'b0;
    assign data[10711] = 16'b0;
    assign data[10712] = ~16'b0;
    assign data[10713] = ~16'b0;
    assign data[10714] = ~16'b0;
    assign data[10715] = ~16'b0;
    assign data[10716] = ~16'b0;
    assign data[10717] = ~16'b0;
    assign data[10718] = ~16'b0;
    assign data[10719] = ~16'b0;
    assign data[10720] = 16'b0;
    assign data[10721] = 16'b0;
    assign data[10722] = ~16'b0;
    assign data[10723] = ~16'b0;
    assign data[10724] = ~16'b0;
    assign data[10725] = ~16'b0;
    assign data[10726] = ~16'b0;
    assign data[10727] = ~16'b0;
    assign data[10728] = ~16'b0;
    assign data[10729] = ~16'b0;
    assign data[10730] = 16'b0;
    assign data[10731] = 16'b0;
    assign data[10732] = ~16'b0;
    assign data[10733] = ~16'b0;
    assign data[10734] = ~16'b0;
    assign data[10735] = ~16'b0;
    assign data[10736] = ~16'b0;
    assign data[10737] = ~16'b0;
    assign data[10738] = ~16'b0;
    assign data[10739] = ~16'b0;
    assign data[10740] = 16'b0;
    assign data[10741] = 16'b0;
    assign data[10742] = ~16'b0;
    assign data[10743] = ~16'b0;
    assign data[10744] = ~16'b0;
    assign data[10745] = ~16'b0;
    assign data[10746] = ~16'b0;
    assign data[10747] = ~16'b0;
    assign data[10748] = ~16'b0;
    assign data[10749] = ~16'b0;
    assign data[10750] = 16'b0;
    assign data[10751] = 16'b0;
    assign data[10752] = ~16'b0;
    assign data[10753] = ~16'b0;
    assign data[10754] = ~16'b0;
    assign data[10755] = ~16'b0;
    assign data[10756] = ~16'b0;
    assign data[10757] = ~16'b0;
    assign data[10758] = ~16'b0;
    assign data[10759] = ~16'b0;
    assign data[10760] = 16'b0;
    assign data[10761] = 16'b0;
    assign data[10762] = ~16'b0;
    assign data[10763] = ~16'b0;
    assign data[10764] = ~16'b0;
    assign data[10765] = ~16'b0;
    assign data[10766] = ~16'b0;
    assign data[10767] = ~16'b0;
    assign data[10768] = ~16'b0;
    assign data[10769] = ~16'b0;
    assign data[10770] = 16'b0;
    assign data[10771] = 16'b0;
    assign data[10772] = ~16'b0;
    assign data[10773] = ~16'b0;
    assign data[10774] = ~16'b0;
    assign data[10775] = ~16'b0;
    assign data[10776] = ~16'b0;
    assign data[10777] = ~16'b0;
    assign data[10778] = ~16'b0;
    assign data[10779] = ~16'b0;
    assign data[10780] = 16'b0;
    assign data[10781] = 16'b0;
    assign data[10782] = ~16'b0;
    assign data[10783] = ~16'b0;
    assign data[10784] = ~16'b0;
    assign data[10785] = ~16'b0;
    assign data[10786] = ~16'b0;
    assign data[10787] = ~16'b0;
    assign data[10788] = ~16'b0;
    assign data[10789] = ~16'b0;
    assign data[10790] = 16'b0;
    assign data[10791] = 16'b0;
    assign data[10792] = ~16'b0;
    assign data[10793] = ~16'b0;
    assign data[10794] = ~16'b0;
    assign data[10795] = ~16'b0;
    assign data[10796] = ~16'b0;
    assign data[10797] = ~16'b0;
    assign data[10798] = ~16'b0;
    assign data[10799] = ~16'b0;
    assign data[10800] = 16'b0;
    assign data[10801] = 16'b0;
    assign data[10802] = ~16'b0;
    assign data[10803] = ~16'b0;
    assign data[10804] = ~16'b0;
    assign data[10805] = ~16'b0;
    assign data[10806] = ~16'b0;
    assign data[10807] = ~16'b0;
    assign data[10808] = ~16'b0;
    assign data[10809] = ~16'b0;
    assign data[10810] = 16'b0;
    assign data[10811] = 16'b0;
    assign data[10812] = ~16'b0;
    assign data[10813] = ~16'b0;
    assign data[10814] = ~16'b0;
    assign data[10815] = ~16'b0;
    assign data[10816] = ~16'b0;
    assign data[10817] = ~16'b0;
    assign data[10818] = ~16'b0;
    assign data[10819] = ~16'b0;
    assign data[10820] = 16'b0;
    assign data[10821] = 16'b0;
    assign data[10822] = ~16'b0;
    assign data[10823] = ~16'b0;
    assign data[10824] = ~16'b0;
    assign data[10825] = ~16'b0;
    assign data[10826] = ~16'b0;
    assign data[10827] = ~16'b0;
    assign data[10828] = ~16'b0;
    assign data[10829] = ~16'b0;
    assign data[10830] = 16'b0;
    assign data[10831] = 16'b0;
    assign data[10832] = ~16'b0;
    assign data[10833] = ~16'b0;
    assign data[10834] = ~16'b0;
    assign data[10835] = ~16'b0;
    assign data[10836] = ~16'b0;
    assign data[10837] = ~16'b0;
    assign data[10838] = ~16'b0;
    assign data[10839] = ~16'b0;
    assign data[10840] = 16'b0;
    assign data[10841] = 16'b0;
    assign data[10842] = ~16'b0;
    assign data[10843] = ~16'b0;
    assign data[10844] = ~16'b0;
    assign data[10845] = ~16'b0;
    assign data[10846] = ~16'b0;
    assign data[10847] = ~16'b0;
    assign data[10848] = ~16'b0;
    assign data[10849] = ~16'b0;
    assign data[10850] = 16'b0;
    assign data[10851] = 16'b0;
    assign data[10852] = 16'b0;
    assign data[10853] = 16'b0;
    assign data[10854] = 16'b0;
    assign data[10855] = 16'b0;
    assign data[10856] = 16'b0;
    assign data[10857] = 16'b0;
    assign data[10858] = 16'b0;
    assign data[10859] = 16'b0;
    assign data[10860] = 16'b0;
    assign data[10861] = 16'b0;
    assign data[10862] = 16'b0;
    assign data[10863] = 16'b0;
    assign data[10864] = 16'b0;
    assign data[10865] = 16'b0;
    assign data[10866] = 16'b0;
    assign data[10867] = 16'b0;
    assign data[10868] = 16'b0;
    assign data[10869] = 16'b0;
    assign data[10870] = ~16'b0;
    assign data[10871] = ~16'b0;
    assign data[10872] = ~16'b0;
    assign data[10873] = ~16'b0;
    assign data[10874] = ~16'b0;
    assign data[10875] = ~16'b0;
    assign data[10876] = ~16'b0;
    assign data[10877] = ~16'b0;
    assign data[10878] = ~16'b0;
    assign data[10879] = ~16'b0;
    assign data[10880] = ~16'b0;
    assign data[10881] = ~16'b0;
    assign data[10882] = ~16'b0;
    assign data[10883] = ~16'b0;
    assign data[10884] = ~16'b0;
    assign data[10885] = ~16'b0;
    assign data[10886] = ~16'b0;
    assign data[10887] = ~16'b0;
    assign data[10888] = ~16'b0;
    assign data[10889] = ~16'b0;
    assign data[10890] = ~16'b0;
    assign data[10891] = ~16'b0;
    assign data[10892] = ~16'b0;
    assign data[10893] = ~16'b0;
    assign data[10894] = ~16'b0;
    assign data[10895] = ~16'b0;
    assign data[10896] = ~16'b0;
    assign data[10897] = ~16'b0;
    assign data[10898] = ~16'b0;
    assign data[10899] = ~16'b0;
    assign data[10900] = ~16'b0;
    assign data[10901] = ~16'b0;
    assign data[10902] = ~16'b0;
    assign data[10903] = ~16'b0;
    assign data[10904] = ~16'b0;
    assign data[10905] = ~16'b0;
    assign data[10906] = ~16'b0;
    assign data[10907] = ~16'b0;
    assign data[10908] = ~16'b0;
    assign data[10909] = ~16'b0;
    assign data[10910] = ~16'b0;
    assign data[10911] = ~16'b0;
    assign data[10912] = ~16'b0;
    assign data[10913] = ~16'b0;
    assign data[10914] = ~16'b0;
    assign data[10915] = ~16'b0;
    assign data[10916] = ~16'b0;
    assign data[10917] = ~16'b0;
    assign data[10918] = ~16'b0;
    assign data[10919] = ~16'b0;
    assign data[10920] = ~16'b0;
    assign data[10921] = ~16'b0;
    assign data[10922] = ~16'b0;
    assign data[10923] = ~16'b0;
    assign data[10924] = ~16'b0;
    assign data[10925] = ~16'b0;
    assign data[10926] = ~16'b0;
    assign data[10927] = ~16'b0;
    assign data[10928] = ~16'b0;
    assign data[10929] = ~16'b0;
    assign data[10930] = ~16'b0;
    assign data[10931] = ~16'b0;
    assign data[10932] = ~16'b0;
    assign data[10933] = ~16'b0;
    assign data[10934] = ~16'b0;
    assign data[10935] = ~16'b0;
    assign data[10936] = ~16'b0;
    assign data[10937] = ~16'b0;
    assign data[10938] = ~16'b0;
    assign data[10939] = ~16'b0;
    assign data[10940] = ~16'b0;
    assign data[10941] = ~16'b0;
    assign data[10942] = ~16'b0;
    assign data[10943] = ~16'b0;
    assign data[10944] = ~16'b0;
    assign data[10945] = ~16'b0;
    assign data[10946] = ~16'b0;
    assign data[10947] = ~16'b0;
    assign data[10948] = ~16'b0;
    assign data[10949] = ~16'b0;
    assign data[10950] = ~16'b0;
    assign data[10951] = ~16'b0;
    assign data[10952] = ~16'b0;
    assign data[10953] = ~16'b0;
    assign data[10954] = ~16'b0;
    assign data[10955] = ~16'b0;
    assign data[10956] = ~16'b0;
    assign data[10957] = ~16'b0;
    assign data[10958] = ~16'b0;
    assign data[10959] = ~16'b0;
    assign data[10960] = ~16'b0;
    assign data[10961] = ~16'b0;
    assign data[10962] = ~16'b0;
    assign data[10963] = ~16'b0;
    assign data[10964] = ~16'b0;
    assign data[10965] = ~16'b0;
    assign data[10966] = ~16'b0;
    assign data[10967] = ~16'b0;
    assign data[10968] = ~16'b0;
    assign data[10969] = ~16'b0;
    assign data[10970] = ~16'b0;
    assign data[10971] = ~16'b0;
    assign data[10972] = ~16'b0;
    assign data[10973] = ~16'b0;
    assign data[10974] = ~16'b0;
    assign data[10975] = ~16'b0;
    assign data[10976] = ~16'b0;
    assign data[10977] = ~16'b0;
    assign data[10978] = ~16'b0;
    assign data[10979] = ~16'b0;
    assign data[10980] = ~16'b0;
    assign data[10981] = ~16'b0;
    assign data[10982] = ~16'b0;
    assign data[10983] = ~16'b0;
    assign data[10984] = ~16'b0;
    assign data[10985] = ~16'b0;
    assign data[10986] = ~16'b0;
    assign data[10987] = ~16'b0;
    assign data[10988] = ~16'b0;
    assign data[10989] = ~16'b0;
    assign data[10990] = ~16'b0;
    assign data[10991] = ~16'b0;
    assign data[10992] = ~16'b0;
    assign data[10993] = ~16'b0;
    assign data[10994] = ~16'b0;
    assign data[10995] = ~16'b0;
    assign data[10996] = ~16'b0;
    assign data[10997] = ~16'b0;
    assign data[10998] = ~16'b0;
    assign data[10999] = ~16'b0;
    assign data[11000] = ~16'b0;
    assign data[11001] = ~16'b0;
    assign data[11002] = ~16'b0;
    assign data[11003] = ~16'b0;
    assign data[11004] = ~16'b0;
    assign data[11005] = ~16'b0;
    assign data[11006] = ~16'b0;
    assign data[11007] = ~16'b0;
    assign data[11008] = ~16'b0;
    assign data[11009] = ~16'b0;
    assign data[11010] = ~16'b0;
    assign data[11011] = ~16'b0;
    assign data[11012] = ~16'b0;
    assign data[11013] = ~16'b0;
    assign data[11014] = ~16'b0;
    assign data[11015] = ~16'b0;
    assign data[11016] = ~16'b0;
    assign data[11017] = ~16'b0;
    assign data[11018] = ~16'b0;
    assign data[11019] = ~16'b0;
    assign data[11020] = ~16'b0;
    assign data[11021] = ~16'b0;
    assign data[11022] = ~16'b0;
    assign data[11023] = ~16'b0;
    assign data[11024] = ~16'b0;
    assign data[11025] = ~16'b0;
    assign data[11026] = ~16'b0;
    assign data[11027] = ~16'b0;
    assign data[11028] = ~16'b0;
    assign data[11029] = ~16'b0;
    assign data[11030] = ~16'b0;
    assign data[11031] = ~16'b0;
    assign data[11032] = ~16'b0;
    assign data[11033] = ~16'b0;
    assign data[11034] = ~16'b0;
    assign data[11035] = ~16'b0;
    assign data[11036] = ~16'b0;
    assign data[11037] = ~16'b0;
    assign data[11038] = ~16'b0;
    assign data[11039] = ~16'b0;
    assign data[11040] = ~16'b0;
    assign data[11041] = ~16'b0;
    assign data[11042] = ~16'b0;
    assign data[11043] = ~16'b0;
    assign data[11044] = ~16'b0;
    assign data[11045] = ~16'b0;
    assign data[11046] = ~16'b0;
    assign data[11047] = ~16'b0;
    assign data[11048] = ~16'b0;
    assign data[11049] = ~16'b0;
    assign data[11050] = ~16'b0;
    assign data[11051] = ~16'b0;
    assign data[11052] = ~16'b0;
    assign data[11053] = ~16'b0;
    assign data[11054] = ~16'b0;
    assign data[11055] = ~16'b0;
    assign data[11056] = ~16'b0;
    assign data[11057] = ~16'b0;
    assign data[11058] = ~16'b0;
    assign data[11059] = ~16'b0;
    assign data[11060] = ~16'b0;
    assign data[11061] = ~16'b0;
    assign data[11062] = ~16'b0;
    assign data[11063] = ~16'b0;
    assign data[11064] = ~16'b0;
    assign data[11065] = ~16'b0;
    assign data[11066] = ~16'b0;
    assign data[11067] = ~16'b0;
    assign data[11068] = ~16'b0;
    assign data[11069] = ~16'b0;
    assign data[11070] = 16'b0;
    assign data[11071] = 16'b0;
    assign data[11072] = 16'b0;
    assign data[11073] = 16'b0;
    assign data[11074] = 16'b0;
    assign data[11075] = 16'b0;
    assign data[11076] = 16'b0;
    assign data[11077] = 16'b0;
    assign data[11078] = 16'b0;
    assign data[11079] = 16'b0;
    assign data[11080] = 16'b0;
    assign data[11081] = 16'b0;
    assign data[11082] = 16'b0;
    assign data[11083] = 16'b0;
    assign data[11084] = 16'b0;
    assign data[11085] = 16'b0;
    assign data[11086] = 16'b0;
    assign data[11087] = 16'b0;
    assign data[11088] = 16'b0;
    assign data[11089] = 16'b0;
    assign data[11090] = 16'b0;
    assign data[11091] = 16'b0;
    assign data[11092] = ~16'b0;
    assign data[11093] = ~16'b0;
    assign data[11094] = ~16'b0;
    assign data[11095] = ~16'b0;
    assign data[11096] = ~16'b0;
    assign data[11097] = ~16'b0;
    assign data[11098] = ~16'b0;
    assign data[11099] = ~16'b0;
    assign data[11100] = 16'b0;
    assign data[11101] = 16'b0;
    assign data[11102] = ~16'b0;
    assign data[11103] = ~16'b0;
    assign data[11104] = ~16'b0;
    assign data[11105] = ~16'b0;
    assign data[11106] = ~16'b0;
    assign data[11107] = ~16'b0;
    assign data[11108] = ~16'b0;
    assign data[11109] = ~16'b0;
    assign data[11110] = 16'b0;
    assign data[11111] = 16'b0;
    assign data[11112] = ~16'b0;
    assign data[11113] = ~16'b0;
    assign data[11114] = ~16'b0;
    assign data[11115] = ~16'b0;
    assign data[11116] = ~16'b0;
    assign data[11117] = ~16'b0;
    assign data[11118] = ~16'b0;
    assign data[11119] = ~16'b0;
    assign data[11120] = 16'b0;
    assign data[11121] = 16'b0;
    assign data[11122] = ~16'b0;
    assign data[11123] = ~16'b0;
    assign data[11124] = ~16'b0;
    assign data[11125] = ~16'b0;
    assign data[11126] = ~16'b0;
    assign data[11127] = ~16'b0;
    assign data[11128] = ~16'b0;
    assign data[11129] = ~16'b0;
    assign data[11130] = 16'b0;
    assign data[11131] = 16'b0;
    assign data[11132] = ~16'b0;
    assign data[11133] = ~16'b0;
    assign data[11134] = ~16'b0;
    assign data[11135] = ~16'b0;
    assign data[11136] = ~16'b0;
    assign data[11137] = ~16'b0;
    assign data[11138] = ~16'b0;
    assign data[11139] = ~16'b0;
    assign data[11140] = 16'b0;
    assign data[11141] = 16'b0;
    assign data[11142] = ~16'b0;
    assign data[11143] = ~16'b0;
    assign data[11144] = ~16'b0;
    assign data[11145] = ~16'b0;
    assign data[11146] = ~16'b0;
    assign data[11147] = ~16'b0;
    assign data[11148] = ~16'b0;
    assign data[11149] = ~16'b0;
    assign data[11150] = 16'b0;
    assign data[11151] = 16'b0;
    assign data[11152] = ~16'b0;
    assign data[11153] = ~16'b0;
    assign data[11154] = ~16'b0;
    assign data[11155] = ~16'b0;
    assign data[11156] = ~16'b0;
    assign data[11157] = ~16'b0;
    assign data[11158] = ~16'b0;
    assign data[11159] = ~16'b0;
    assign data[11160] = 16'b0;
    assign data[11161] = 16'b0;
    assign data[11162] = ~16'b0;
    assign data[11163] = ~16'b0;
    assign data[11164] = ~16'b0;
    assign data[11165] = ~16'b0;
    assign data[11166] = ~16'b0;
    assign data[11167] = ~16'b0;
    assign data[11168] = ~16'b0;
    assign data[11169] = ~16'b0;
    assign data[11170] = 16'b0;
    assign data[11171] = 16'b0;
    assign data[11172] = ~16'b0;
    assign data[11173] = ~16'b0;
    assign data[11174] = ~16'b0;
    assign data[11175] = ~16'b0;
    assign data[11176] = ~16'b0;
    assign data[11177] = ~16'b0;
    assign data[11178] = ~16'b0;
    assign data[11179] = ~16'b0;
    assign data[11180] = 16'b0;
    assign data[11181] = 16'b0;
    assign data[11182] = ~16'b0;
    assign data[11183] = ~16'b0;
    assign data[11184] = ~16'b0;
    assign data[11185] = ~16'b0;
    assign data[11186] = ~16'b0;
    assign data[11187] = ~16'b0;
    assign data[11188] = ~16'b0;
    assign data[11189] = ~16'b0;
    assign data[11190] = 16'b0;
    assign data[11191] = 16'b0;
    assign data[11192] = ~16'b0;
    assign data[11193] = ~16'b0;
    assign data[11194] = ~16'b0;
    assign data[11195] = ~16'b0;
    assign data[11196] = ~16'b0;
    assign data[11197] = ~16'b0;
    assign data[11198] = ~16'b0;
    assign data[11199] = ~16'b0;
    assign data[11200] = 16'b0;
    assign data[11201] = 16'b0;
    assign data[11202] = ~16'b0;
    assign data[11203] = ~16'b0;
    assign data[11204] = ~16'b0;
    assign data[11205] = ~16'b0;
    assign data[11206] = ~16'b0;
    assign data[11207] = ~16'b0;
    assign data[11208] = ~16'b0;
    assign data[11209] = ~16'b0;
    assign data[11210] = 16'b0;
    assign data[11211] = 16'b0;
    assign data[11212] = ~16'b0;
    assign data[11213] = ~16'b0;
    assign data[11214] = ~16'b0;
    assign data[11215] = ~16'b0;
    assign data[11216] = ~16'b0;
    assign data[11217] = ~16'b0;
    assign data[11218] = ~16'b0;
    assign data[11219] = ~16'b0;
    assign data[11220] = 16'b0;
    assign data[11221] = 16'b0;
    assign data[11222] = ~16'b0;
    assign data[11223] = ~16'b0;
    assign data[11224] = ~16'b0;
    assign data[11225] = ~16'b0;
    assign data[11226] = ~16'b0;
    assign data[11227] = ~16'b0;
    assign data[11228] = ~16'b0;
    assign data[11229] = ~16'b0;
    assign data[11230] = 16'b0;
    assign data[11231] = 16'b0;
    assign data[11232] = ~16'b0;
    assign data[11233] = ~16'b0;
    assign data[11234] = ~16'b0;
    assign data[11235] = ~16'b0;
    assign data[11236] = ~16'b0;
    assign data[11237] = ~16'b0;
    assign data[11238] = ~16'b0;
    assign data[11239] = ~16'b0;
    assign data[11240] = 16'b0;
    assign data[11241] = 16'b0;
    assign data[11242] = ~16'b0;
    assign data[11243] = ~16'b0;
    assign data[11244] = ~16'b0;
    assign data[11245] = ~16'b0;
    assign data[11246] = ~16'b0;
    assign data[11247] = ~16'b0;
    assign data[11248] = ~16'b0;
    assign data[11249] = ~16'b0;
    assign data[11250] = 16'b0;
    assign data[11251] = 16'b0;
    assign data[11252] = ~16'b0;
    assign data[11253] = ~16'b0;
    assign data[11254] = ~16'b0;
    assign data[11255] = ~16'b0;
    assign data[11256] = ~16'b0;
    assign data[11257] = ~16'b0;
    assign data[11258] = ~16'b0;
    assign data[11259] = ~16'b0;
    assign data[11260] = 16'b0;
    assign data[11261] = 16'b0;
    assign data[11262] = ~16'b0;
    assign data[11263] = ~16'b0;
    assign data[11264] = ~16'b0;
    assign data[11265] = ~16'b0;
    assign data[11266] = ~16'b0;
    assign data[11267] = ~16'b0;
    assign data[11268] = ~16'b0;
    assign data[11269] = ~16'b0;
    assign data[11270] = 16'b0;
    assign data[11271] = 16'b0;
    assign data[11272] = 16'b0;
    assign data[11273] = 16'b0;
    assign data[11274] = 16'b0;
    assign data[11275] = 16'b0;
    assign data[11276] = 16'b0;
    assign data[11277] = 16'b0;
    assign data[11278] = 16'b0;
    assign data[11279] = 16'b0;
    assign data[11280] = 16'b0;
    assign data[11281] = 16'b0;
    assign data[11282] = 16'b0;
    assign data[11283] = 16'b0;
    assign data[11284] = 16'b0;
    assign data[11285] = 16'b0;
    assign data[11286] = 16'b0;
    assign data[11287] = 16'b0;
    assign data[11288] = 16'b0;
    assign data[11289] = 16'b0;
    assign data[11290] = ~16'b0;
    assign data[11291] = ~16'b0;
    assign data[11292] = ~16'b0;
    assign data[11293] = ~16'b0;
    assign data[11294] = ~16'b0;
    assign data[11295] = ~16'b0;
    assign data[11296] = ~16'b0;
    assign data[11297] = ~16'b0;
    assign data[11298] = ~16'b0;
    assign data[11299] = ~16'b0;
    assign data[11300] = ~16'b0;
    assign data[11301] = ~16'b0;
    assign data[11302] = ~16'b0;
    assign data[11303] = ~16'b0;
    assign data[11304] = ~16'b0;
    assign data[11305] = ~16'b0;
    assign data[11306] = ~16'b0;
    assign data[11307] = ~16'b0;
    assign data[11308] = ~16'b0;
    assign data[11309] = ~16'b0;
    assign data[11310] = ~16'b0;
    assign data[11311] = ~16'b0;
    assign data[11312] = ~16'b0;
    assign data[11313] = ~16'b0;
    assign data[11314] = ~16'b0;
    assign data[11315] = ~16'b0;
    assign data[11316] = ~16'b0;
    assign data[11317] = ~16'b0;
    assign data[11318] = ~16'b0;
    assign data[11319] = ~16'b0;
    assign data[11320] = ~16'b0;
    assign data[11321] = ~16'b0;
    assign data[11322] = ~16'b0;
    assign data[11323] = ~16'b0;
    assign data[11324] = ~16'b0;
    assign data[11325] = ~16'b0;
    assign data[11326] = ~16'b0;
    assign data[11327] = ~16'b0;
    assign data[11328] = ~16'b0;
    assign data[11329] = ~16'b0;
    assign data[11330] = ~16'b0;
    assign data[11331] = ~16'b0;
    assign data[11332] = ~16'b0;
    assign data[11333] = ~16'b0;
    assign data[11334] = ~16'b0;
    assign data[11335] = ~16'b0;
    assign data[11336] = ~16'b0;
    assign data[11337] = ~16'b0;
    assign data[11338] = ~16'b0;
    assign data[11339] = ~16'b0;
    assign data[11340] = ~16'b0;
    assign data[11341] = ~16'b0;
    assign data[11342] = ~16'b0;
    assign data[11343] = ~16'b0;
    assign data[11344] = ~16'b0;
    assign data[11345] = ~16'b0;
    assign data[11346] = ~16'b0;
    assign data[11347] = ~16'b0;
    assign data[11348] = ~16'b0;
    assign data[11349] = ~16'b0;
    assign data[11350] = ~16'b0;
    assign data[11351] = ~16'b0;
    assign data[11352] = ~16'b0;
    assign data[11353] = ~16'b0;
    assign data[11354] = ~16'b0;
    assign data[11355] = ~16'b0;
    assign data[11356] = ~16'b0;
    assign data[11357] = ~16'b0;
    assign data[11358] = ~16'b0;
    assign data[11359] = ~16'b0;
    assign data[11360] = ~16'b0;
    assign data[11361] = ~16'b0;
    assign data[11362] = ~16'b0;
    assign data[11363] = ~16'b0;
    assign data[11364] = ~16'b0;
    assign data[11365] = ~16'b0;
    assign data[11366] = ~16'b0;
    assign data[11367] = ~16'b0;
    assign data[11368] = ~16'b0;
    assign data[11369] = ~16'b0;
    assign data[11370] = ~16'b0;
    assign data[11371] = ~16'b0;
    assign data[11372] = ~16'b0;
    assign data[11373] = ~16'b0;
    assign data[11374] = ~16'b0;
    assign data[11375] = ~16'b0;
    assign data[11376] = ~16'b0;
    assign data[11377] = ~16'b0;
    assign data[11378] = ~16'b0;
    assign data[11379] = ~16'b0;
    assign data[11380] = ~16'b0;
    assign data[11381] = ~16'b0;
    assign data[11382] = ~16'b0;
    assign data[11383] = ~16'b0;
    assign data[11384] = ~16'b0;
    assign data[11385] = ~16'b0;
    assign data[11386] = ~16'b0;
    assign data[11387] = ~16'b0;
    assign data[11388] = ~16'b0;
    assign data[11389] = ~16'b0;
    assign data[11390] = ~16'b0;
    assign data[11391] = ~16'b0;
    assign data[11392] = ~16'b0;
    assign data[11393] = ~16'b0;
    assign data[11394] = ~16'b0;
    assign data[11395] = ~16'b0;
    assign data[11396] = ~16'b0;
    assign data[11397] = ~16'b0;
    assign data[11398] = ~16'b0;
    assign data[11399] = ~16'b0;
    assign data[11400] = ~16'b0;
    assign data[11401] = ~16'b0;
    assign data[11402] = ~16'b0;
    assign data[11403] = ~16'b0;
    assign data[11404] = ~16'b0;
    assign data[11405] = ~16'b0;
    assign data[11406] = ~16'b0;
    assign data[11407] = ~16'b0;
    assign data[11408] = ~16'b0;
    assign data[11409] = ~16'b0;
    assign data[11410] = ~16'b0;
    assign data[11411] = ~16'b0;
    assign data[11412] = ~16'b0;
    assign data[11413] = ~16'b0;
    assign data[11414] = ~16'b0;
    assign data[11415] = ~16'b0;
    assign data[11416] = ~16'b0;
    assign data[11417] = ~16'b0;
    assign data[11418] = ~16'b0;
    assign data[11419] = ~16'b0;
    assign data[11420] = ~16'b0;
    assign data[11421] = ~16'b0;
    assign data[11422] = ~16'b0;
    assign data[11423] = ~16'b0;
    assign data[11424] = ~16'b0;
    assign data[11425] = ~16'b0;
    assign data[11426] = ~16'b0;
    assign data[11427] = ~16'b0;
    assign data[11428] = ~16'b0;
    assign data[11429] = ~16'b0;
    assign data[11430] = 16'b0;
    assign data[11431] = 16'b0;
    assign data[11432] = 16'b0;
    assign data[11433] = 16'b0;
    assign data[11434] = 16'b0;
    assign data[11435] = 16'b0;
    assign data[11436] = 16'b0;
    assign data[11437] = 16'b0;
    assign data[11438] = 16'b0;
    assign data[11439] = 16'b0;
    assign data[11440] = 16'b0;
    assign data[11441] = 16'b0;
    assign data[11442] = 16'b0;
    assign data[11443] = 16'b0;
    assign data[11444] = 16'b0;
    assign data[11445] = 16'b0;
    assign data[11446] = 16'b0;
    assign data[11447] = 16'b0;
    assign data[11448] = 16'b0;
    assign data[11449] = 16'b0;
    assign data[11450] = 16'b0;
    assign data[11451] = 16'b0;
    assign data[11452] = ~16'b0;
    assign data[11453] = ~16'b0;
    assign data[11454] = ~16'b0;
    assign data[11455] = ~16'b0;
    assign data[11456] = ~16'b0;
    assign data[11457] = ~16'b0;
    assign data[11458] = ~16'b0;
    assign data[11459] = ~16'b0;
    assign data[11460] = 16'b0;
    assign data[11461] = 16'b0;
    assign data[11462] = ~16'b0;
    assign data[11463] = ~16'b0;
    assign data[11464] = ~16'b0;
    assign data[11465] = ~16'b0;
    assign data[11466] = ~16'b0;
    assign data[11467] = ~16'b0;
    assign data[11468] = ~16'b0;
    assign data[11469] = ~16'b0;
    assign data[11470] = 16'b0;
    assign data[11471] = 16'b0;
    assign data[11472] = ~16'b0;
    assign data[11473] = ~16'b0;
    assign data[11474] = ~16'b0;
    assign data[11475] = ~16'b0;
    assign data[11476] = ~16'b0;
    assign data[11477] = ~16'b0;
    assign data[11478] = ~16'b0;
    assign data[11479] = ~16'b0;
    assign data[11480] = 16'b0;
    assign data[11481] = 16'b0;
    assign data[11482] = ~16'b0;
    assign data[11483] = ~16'b0;
    assign data[11484] = ~16'b0;
    assign data[11485] = ~16'b0;
    assign data[11486] = ~16'b0;
    assign data[11487] = ~16'b0;
    assign data[11488] = ~16'b0;
    assign data[11489] = ~16'b0;
    assign data[11490] = 16'b0;
    assign data[11491] = 16'b0;
    assign data[11492] = ~16'b0;
    assign data[11493] = ~16'b0;
    assign data[11494] = ~16'b0;
    assign data[11495] = ~16'b0;
    assign data[11496] = ~16'b0;
    assign data[11497] = ~16'b0;
    assign data[11498] = ~16'b0;
    assign data[11499] = ~16'b0;
    assign data[11500] = 16'b0;
    assign data[11501] = 16'b0;
    assign data[11502] = ~16'b0;
    assign data[11503] = ~16'b0;
    assign data[11504] = ~16'b0;
    assign data[11505] = ~16'b0;
    assign data[11506] = ~16'b0;
    assign data[11507] = ~16'b0;
    assign data[11508] = ~16'b0;
    assign data[11509] = ~16'b0;
    assign data[11510] = 16'b0;
    assign data[11511] = 16'b0;
    assign data[11512] = ~16'b0;
    assign data[11513] = ~16'b0;
    assign data[11514] = ~16'b0;
    assign data[11515] = ~16'b0;
    assign data[11516] = ~16'b0;
    assign data[11517] = ~16'b0;
    assign data[11518] = ~16'b0;
    assign data[11519] = ~16'b0;
    assign data[11520] = 16'b0;
    assign data[11521] = 16'b0;
    assign data[11522] = ~16'b0;
    assign data[11523] = ~16'b0;
    assign data[11524] = ~16'b0;
    assign data[11525] = ~16'b0;
    assign data[11526] = ~16'b0;
    assign data[11527] = ~16'b0;
    assign data[11528] = ~16'b0;
    assign data[11529] = ~16'b0;
    assign data[11530] = 16'b0;
    assign data[11531] = 16'b0;
    assign data[11532] = ~16'b0;
    assign data[11533] = ~16'b0;
    assign data[11534] = ~16'b0;
    assign data[11535] = ~16'b0;
    assign data[11536] = ~16'b0;
    assign data[11537] = ~16'b0;
    assign data[11538] = ~16'b0;
    assign data[11539] = ~16'b0;
    assign data[11540] = 16'b0;
    assign data[11541] = 16'b0;
    assign data[11542] = ~16'b0;
    assign data[11543] = ~16'b0;
    assign data[11544] = ~16'b0;
    assign data[11545] = ~16'b0;
    assign data[11546] = ~16'b0;
    assign data[11547] = ~16'b0;
    assign data[11548] = ~16'b0;
    assign data[11549] = ~16'b0;
    assign data[11550] = 16'b0;
    assign data[11551] = 16'b0;
    assign data[11552] = ~16'b0;
    assign data[11553] = ~16'b0;
    assign data[11554] = ~16'b0;
    assign data[11555] = ~16'b0;
    assign data[11556] = ~16'b0;
    assign data[11557] = ~16'b0;
    assign data[11558] = ~16'b0;
    assign data[11559] = ~16'b0;
    assign data[11560] = 16'b0;
    assign data[11561] = 16'b0;
    assign data[11562] = ~16'b0;
    assign data[11563] = ~16'b0;
    assign data[11564] = ~16'b0;
    assign data[11565] = ~16'b0;
    assign data[11566] = ~16'b0;
    assign data[11567] = ~16'b0;
    assign data[11568] = ~16'b0;
    assign data[11569] = ~16'b0;
    assign data[11570] = 16'b0;
    assign data[11571] = 16'b0;
    assign data[11572] = ~16'b0;
    assign data[11573] = ~16'b0;
    assign data[11574] = ~16'b0;
    assign data[11575] = ~16'b0;
    assign data[11576] = ~16'b0;
    assign data[11577] = ~16'b0;
    assign data[11578] = ~16'b0;
    assign data[11579] = ~16'b0;
    assign data[11580] = 16'b0;
    assign data[11581] = 16'b0;
    assign data[11582] = ~16'b0;
    assign data[11583] = ~16'b0;
    assign data[11584] = ~16'b0;
    assign data[11585] = ~16'b0;
    assign data[11586] = ~16'b0;
    assign data[11587] = ~16'b0;
    assign data[11588] = ~16'b0;
    assign data[11589] = ~16'b0;
    assign data[11590] = 16'b0;
    assign data[11591] = 16'b0;
    assign data[11592] = ~16'b0;
    assign data[11593] = ~16'b0;
    assign data[11594] = ~16'b0;
    assign data[11595] = ~16'b0;
    assign data[11596] = ~16'b0;
    assign data[11597] = ~16'b0;
    assign data[11598] = ~16'b0;
    assign data[11599] = ~16'b0;
    assign data[11600] = 16'b0;
    assign data[11601] = 16'b0;
    assign data[11602] = ~16'b0;
    assign data[11603] = ~16'b0;
    assign data[11604] = ~16'b0;
    assign data[11605] = ~16'b0;
    assign data[11606] = ~16'b0;
    assign data[11607] = ~16'b0;
    assign data[11608] = ~16'b0;
    assign data[11609] = ~16'b0;
    assign data[11610] = 16'b0;
    assign data[11611] = 16'b0;
    assign data[11612] = ~16'b0;
    assign data[11613] = ~16'b0;
    assign data[11614] = ~16'b0;
    assign data[11615] = ~16'b0;
    assign data[11616] = ~16'b0;
    assign data[11617] = ~16'b0;
    assign data[11618] = ~16'b0;
    assign data[11619] = ~16'b0;
    assign data[11620] = 16'b0;
    assign data[11621] = 16'b0;
    assign data[11622] = ~16'b0;
    assign data[11623] = ~16'b0;
    assign data[11624] = ~16'b0;
    assign data[11625] = ~16'b0;
    assign data[11626] = ~16'b0;
    assign data[11627] = ~16'b0;
    assign data[11628] = ~16'b0;
    assign data[11629] = ~16'b0;
    assign data[11630] = 16'b0;
    assign data[11631] = 16'b0;
    assign data[11632] = ~16'b0;
    assign data[11633] = ~16'b0;
    assign data[11634] = ~16'b0;
    assign data[11635] = ~16'b0;
    assign data[11636] = ~16'b0;
    assign data[11637] = ~16'b0;
    assign data[11638] = ~16'b0;
    assign data[11639] = ~16'b0;
    assign data[11640] = 16'b0;
    assign data[11641] = 16'b0;
    assign data[11642] = ~16'b0;
    assign data[11643] = ~16'b0;
    assign data[11644] = ~16'b0;
    assign data[11645] = ~16'b0;
    assign data[11646] = ~16'b0;
    assign data[11647] = ~16'b0;
    assign data[11648] = ~16'b0;
    assign data[11649] = ~16'b0;
    assign data[11650] = 16'b0;
    assign data[11651] = 16'b0;
    assign data[11652] = ~16'b0;
    assign data[11653] = ~16'b0;
    assign data[11654] = ~16'b0;
    assign data[11655] = ~16'b0;
    assign data[11656] = ~16'b0;
    assign data[11657] = ~16'b0;
    assign data[11658] = ~16'b0;
    assign data[11659] = ~16'b0;
    assign data[11660] = 16'b0;
    assign data[11661] = 16'b0;
    assign data[11662] = ~16'b0;
    assign data[11663] = ~16'b0;
    assign data[11664] = ~16'b0;
    assign data[11665] = ~16'b0;
    assign data[11666] = ~16'b0;
    assign data[11667] = ~16'b0;
    assign data[11668] = ~16'b0;
    assign data[11669] = ~16'b0;
    assign data[11670] = 16'b0;
    assign data[11671] = 16'b0;
    assign data[11672] = ~16'b0;
    assign data[11673] = ~16'b0;
    assign data[11674] = ~16'b0;
    assign data[11675] = ~16'b0;
    assign data[11676] = ~16'b0;
    assign data[11677] = ~16'b0;
    assign data[11678] = ~16'b0;
    assign data[11679] = ~16'b0;
    assign data[11680] = 16'b0;
    assign data[11681] = 16'b0;
    assign data[11682] = ~16'b0;
    assign data[11683] = ~16'b0;
    assign data[11684] = ~16'b0;
    assign data[11685] = ~16'b0;
    assign data[11686] = ~16'b0;
    assign data[11687] = ~16'b0;
    assign data[11688] = ~16'b0;
    assign data[11689] = ~16'b0;
    assign data[11690] = 16'b0;
    assign data[11691] = 16'b0;
    assign data[11692] = ~16'b0;
    assign data[11693] = ~16'b0;
    assign data[11694] = ~16'b0;
    assign data[11695] = ~16'b0;
    assign data[11696] = ~16'b0;
    assign data[11697] = ~16'b0;
    assign data[11698] = ~16'b0;
    assign data[11699] = ~16'b0;
    assign data[11700] = 16'b0;
    assign data[11701] = 16'b0;
    assign data[11702] = ~16'b0;
    assign data[11703] = ~16'b0;
    assign data[11704] = ~16'b0;
    assign data[11705] = ~16'b0;
    assign data[11706] = ~16'b0;
    assign data[11707] = ~16'b0;
    assign data[11708] = ~16'b0;
    assign data[11709] = ~16'b0;
    assign data[11710] = 16'b0;
    assign data[11711] = 16'b0;
    assign data[11712] = ~16'b0;
    assign data[11713] = ~16'b0;
    assign data[11714] = ~16'b0;
    assign data[11715] = ~16'b0;
    assign data[11716] = ~16'b0;
    assign data[11717] = ~16'b0;
    assign data[11718] = ~16'b0;
    assign data[11719] = ~16'b0;
    assign data[11720] = 16'b0;
    assign data[11721] = 16'b0;
    assign data[11722] = ~16'b0;
    assign data[11723] = ~16'b0;
    assign data[11724] = ~16'b0;
    assign data[11725] = ~16'b0;
    assign data[11726] = ~16'b0;
    assign data[11727] = ~16'b0;
    assign data[11728] = ~16'b0;
    assign data[11729] = ~16'b0;
    assign data[11730] = 16'b0;
    assign data[11731] = 16'b0;
    assign data[11732] = ~16'b0;
    assign data[11733] = ~16'b0;
    assign data[11734] = ~16'b0;
    assign data[11735] = ~16'b0;
    assign data[11736] = ~16'b0;
    assign data[11737] = ~16'b0;
    assign data[11738] = ~16'b0;
    assign data[11739] = ~16'b0;
    assign data[11740] = 16'b0;
    assign data[11741] = 16'b0;
    assign data[11742] = ~16'b0;
    assign data[11743] = ~16'b0;
    assign data[11744] = ~16'b0;
    assign data[11745] = ~16'b0;
    assign data[11746] = ~16'b0;
    assign data[11747] = ~16'b0;
    assign data[11748] = ~16'b0;
    assign data[11749] = ~16'b0;
    assign data[11750] = 16'b0;
    assign data[11751] = 16'b0;
    assign data[11752] = ~16'b0;
    assign data[11753] = ~16'b0;
    assign data[11754] = ~16'b0;
    assign data[11755] = ~16'b0;
    assign data[11756] = ~16'b0;
    assign data[11757] = ~16'b0;
    assign data[11758] = ~16'b0;
    assign data[11759] = ~16'b0;
    assign data[11760] = 16'b0;
    assign data[11761] = 16'b0;
    assign data[11762] = ~16'b0;
    assign data[11763] = ~16'b0;
    assign data[11764] = ~16'b0;
    assign data[11765] = ~16'b0;
    assign data[11766] = ~16'b0;
    assign data[11767] = ~16'b0;
    assign data[11768] = ~16'b0;
    assign data[11769] = ~16'b0;
    assign data[11770] = 16'b0;
    assign data[11771] = 16'b0;
    assign data[11772] = ~16'b0;
    assign data[11773] = ~16'b0;
    assign data[11774] = ~16'b0;
    assign data[11775] = ~16'b0;
    assign data[11776] = ~16'b0;
    assign data[11777] = ~16'b0;
    assign data[11778] = ~16'b0;
    assign data[11779] = ~16'b0;
    assign data[11780] = 16'b0;
    assign data[11781] = 16'b0;
    assign data[11782] = ~16'b0;
    assign data[11783] = ~16'b0;
    assign data[11784] = ~16'b0;
    assign data[11785] = ~16'b0;
    assign data[11786] = ~16'b0;
    assign data[11787] = ~16'b0;
    assign data[11788] = ~16'b0;
    assign data[11789] = ~16'b0;
    assign data[11790] = 16'b0;
    assign data[11791] = 16'b0;
    assign data[11792] = ~16'b0;
    assign data[11793] = ~16'b0;
    assign data[11794] = ~16'b0;
    assign data[11795] = ~16'b0;
    assign data[11796] = ~16'b0;
    assign data[11797] = ~16'b0;
    assign data[11798] = ~16'b0;
    assign data[11799] = ~16'b0;
    assign data[11800] = 16'b0;
    assign data[11801] = 16'b0;
    assign data[11802] = ~16'b0;
    assign data[11803] = ~16'b0;
    assign data[11804] = ~16'b0;
    assign data[11805] = ~16'b0;
    assign data[11806] = ~16'b0;
    assign data[11807] = ~16'b0;
    assign data[11808] = ~16'b0;
    assign data[11809] = ~16'b0;
    assign data[11810] = 16'b0;
    assign data[11811] = 16'b0;
    assign data[11812] = 16'b0;
    assign data[11813] = 16'b0;
    assign data[11814] = 16'b0;
    assign data[11815] = 16'b0;
    assign data[11816] = 16'b0;
    assign data[11817] = 16'b0;
    assign data[11818] = 16'b0;
    assign data[11819] = 16'b0;
    assign data[11820] = 16'b0;
    assign data[11821] = 16'b0;
    assign data[11822] = 16'b0;
    assign data[11823] = 16'b0;
    assign data[11824] = 16'b0;
    assign data[11825] = 16'b0;
    assign data[11826] = 16'b0;
    assign data[11827] = 16'b0;
    assign data[11828] = 16'b0;
    assign data[11829] = 16'b0;
    assign data[11830] = ~16'b0;
    assign data[11831] = ~16'b0;
    assign data[11832] = ~16'b0;
    assign data[11833] = ~16'b0;
    assign data[11834] = ~16'b0;
    assign data[11835] = ~16'b0;
    assign data[11836] = ~16'b0;
    assign data[11837] = ~16'b0;
    assign data[11838] = ~16'b0;
    assign data[11839] = ~16'b0;
    assign data[11840] = ~16'b0;
    assign data[11841] = ~16'b0;
    assign data[11842] = ~16'b0;
    assign data[11843] = ~16'b0;
    assign data[11844] = ~16'b0;
    assign data[11845] = ~16'b0;
    assign data[11846] = ~16'b0;
    assign data[11847] = ~16'b0;
    assign data[11848] = ~16'b0;
    assign data[11849] = ~16'b0;
    assign data[11850] = ~16'b0;
    assign data[11851] = ~16'b0;
    assign data[11852] = ~16'b0;
    assign data[11853] = ~16'b0;
    assign data[11854] = ~16'b0;
    assign data[11855] = ~16'b0;
    assign data[11856] = ~16'b0;
    assign data[11857] = ~16'b0;
    assign data[11858] = ~16'b0;
    assign data[11859] = ~16'b0;
    assign data[11860] = ~16'b0;
    assign data[11861] = ~16'b0;
    assign data[11862] = ~16'b0;
    assign data[11863] = ~16'b0;
    assign data[11864] = ~16'b0;
    assign data[11865] = ~16'b0;
    assign data[11866] = ~16'b0;
    assign data[11867] = ~16'b0;
    assign data[11868] = ~16'b0;
    assign data[11869] = ~16'b0;
    assign data[11870] = ~16'b0;
    assign data[11871] = ~16'b0;
    assign data[11872] = ~16'b0;
    assign data[11873] = ~16'b0;
    assign data[11874] = ~16'b0;
    assign data[11875] = ~16'b0;
    assign data[11876] = ~16'b0;
    assign data[11877] = ~16'b0;
    assign data[11878] = ~16'b0;
    assign data[11879] = ~16'b0;
    assign data[11880] = ~16'b0;
    assign data[11881] = ~16'b0;
    assign data[11882] = ~16'b0;
    assign data[11883] = ~16'b0;
    assign data[11884] = ~16'b0;
    assign data[11885] = ~16'b0;
    assign data[11886] = ~16'b0;
    assign data[11887] = ~16'b0;
    assign data[11888] = ~16'b0;
    assign data[11889] = ~16'b0;
    assign data[11890] = ~16'b0;
    assign data[11891] = ~16'b0;
    assign data[11892] = ~16'b0;
    assign data[11893] = ~16'b0;
    assign data[11894] = ~16'b0;
    assign data[11895] = ~16'b0;
    assign data[11896] = ~16'b0;
    assign data[11897] = ~16'b0;
    assign data[11898] = ~16'b0;
    assign data[11899] = ~16'b0;
    assign data[11900] = ~16'b0;
    assign data[11901] = ~16'b0;
    assign data[11902] = ~16'b0;
    assign data[11903] = ~16'b0;
    assign data[11904] = ~16'b0;
    assign data[11905] = ~16'b0;
    assign data[11906] = ~16'b0;
    assign data[11907] = ~16'b0;
    assign data[11908] = ~16'b0;
    assign data[11909] = ~16'b0;
    assign data[11910] = ~16'b0;
    assign data[11911] = ~16'b0;
    assign data[11912] = ~16'b0;
    assign data[11913] = ~16'b0;
    assign data[11914] = ~16'b0;
    assign data[11915] = ~16'b0;
    assign data[11916] = ~16'b0;
    assign data[11917] = ~16'b0;
    assign data[11918] = ~16'b0;
    assign data[11919] = ~16'b0;
    assign data[11920] = ~16'b0;
    assign data[11921] = ~16'b0;
    assign data[11922] = ~16'b0;
    assign data[11923] = ~16'b0;
    assign data[11924] = ~16'b0;
    assign data[11925] = ~16'b0;
    assign data[11926] = ~16'b0;
    assign data[11927] = ~16'b0;
    assign data[11928] = ~16'b0;
    assign data[11929] = ~16'b0;
    assign data[11930] = ~16'b0;
    assign data[11931] = ~16'b0;
    assign data[11932] = ~16'b0;
    assign data[11933] = ~16'b0;
    assign data[11934] = ~16'b0;
    assign data[11935] = ~16'b0;
    assign data[11936] = ~16'b0;
    assign data[11937] = ~16'b0;
    assign data[11938] = ~16'b0;
    assign data[11939] = ~16'b0;
    assign data[11940] = ~16'b0;
    assign data[11941] = ~16'b0;
    assign data[11942] = ~16'b0;
    assign data[11943] = ~16'b0;
    assign data[11944] = ~16'b0;
    assign data[11945] = ~16'b0;
    assign data[11946] = ~16'b0;
    assign data[11947] = ~16'b0;
    assign data[11948] = ~16'b0;
    assign data[11949] = ~16'b0;
    assign data[11950] = ~16'b0;
    assign data[11951] = ~16'b0;
    assign data[11952] = ~16'b0;
    assign data[11953] = ~16'b0;
    assign data[11954] = ~16'b0;
    assign data[11955] = ~16'b0;
    assign data[11956] = ~16'b0;
    assign data[11957] = ~16'b0;
    assign data[11958] = ~16'b0;
    assign data[11959] = ~16'b0;
    assign data[11960] = 16'b0;
    assign data[11961] = 16'b0;
    assign data[11962] = 16'b0;
    assign data[11963] = 16'b0;
    assign data[11964] = 16'b0;
    assign data[11965] = 16'b0;
    assign data[11966] = 16'b0;
    assign data[11967] = 16'b0;
    assign data[11968] = 16'b0;
    assign data[11969] = 16'b0;
    assign data[11970] = 16'b0;
    assign data[11971] = 16'b0;
    assign data[11972] = 16'b0;
    assign data[11973] = 16'b0;
    assign data[11974] = 16'b0;
    assign data[11975] = 16'b0;
    assign data[11976] = 16'b0;
    assign data[11977] = 16'b0;
    assign data[11978] = 16'b0;
    assign data[11979] = 16'b0;
    assign data[11980] = 16'b0;
    assign data[11981] = 16'b0;
    assign data[11982] = ~16'b0;
    assign data[11983] = ~16'b0;
    assign data[11984] = ~16'b0;
    assign data[11985] = ~16'b0;
    assign data[11986] = ~16'b0;
    assign data[11987] = ~16'b0;
    assign data[11988] = ~16'b0;
    assign data[11989] = ~16'b0;
    assign data[11990] = 16'b0;
    assign data[11991] = 16'b0;
    assign data[11992] = ~16'b0;
    assign data[11993] = ~16'b0;
    assign data[11994] = ~16'b0;
    assign data[11995] = ~16'b0;
    assign data[11996] = ~16'b0;
    assign data[11997] = ~16'b0;
    assign data[11998] = ~16'b0;
    assign data[11999] = ~16'b0;
    assign data[12000] = 16'b0;
    assign data[12001] = 16'b0;
    assign data[12002] = ~16'b0;
    assign data[12003] = ~16'b0;
    assign data[12004] = ~16'b0;
    assign data[12005] = ~16'b0;
    assign data[12006] = ~16'b0;
    assign data[12007] = ~16'b0;
    assign data[12008] = ~16'b0;
    assign data[12009] = ~16'b0;
    assign data[12010] = 16'b0;
    assign data[12011] = 16'b0;
    assign data[12012] = ~16'b0;
    assign data[12013] = ~16'b0;
    assign data[12014] = ~16'b0;
    assign data[12015] = ~16'b0;
    assign data[12016] = ~16'b0;
    assign data[12017] = ~16'b0;
    assign data[12018] = ~16'b0;
    assign data[12019] = ~16'b0;
    assign data[12020] = 16'b0;
    assign data[12021] = 16'b0;
    assign data[12022] = ~16'b0;
    assign data[12023] = ~16'b0;
    assign data[12024] = ~16'b0;
    assign data[12025] = ~16'b0;
    assign data[12026] = ~16'b0;
    assign data[12027] = ~16'b0;
    assign data[12028] = ~16'b0;
    assign data[12029] = ~16'b0;
    assign data[12030] = 16'b0;
    assign data[12031] = 16'b0;
    assign data[12032] = ~16'b0;
    assign data[12033] = ~16'b0;
    assign data[12034] = ~16'b0;
    assign data[12035] = ~16'b0;
    assign data[12036] = ~16'b0;
    assign data[12037] = ~16'b0;
    assign data[12038] = ~16'b0;
    assign data[12039] = ~16'b0;
    assign data[12040] = 16'b0;
    assign data[12041] = 16'b0;
    assign data[12042] = ~16'b0;
    assign data[12043] = ~16'b0;
    assign data[12044] = ~16'b0;
    assign data[12045] = ~16'b0;
    assign data[12046] = ~16'b0;
    assign data[12047] = ~16'b0;
    assign data[12048] = ~16'b0;
    assign data[12049] = ~16'b0;
    assign data[12050] = 16'b0;
    assign data[12051] = 16'b0;
    assign data[12052] = ~16'b0;
    assign data[12053] = ~16'b0;
    assign data[12054] = ~16'b0;
    assign data[12055] = ~16'b0;
    assign data[12056] = ~16'b0;
    assign data[12057] = ~16'b0;
    assign data[12058] = ~16'b0;
    assign data[12059] = ~16'b0;
    assign data[12060] = 16'b0;
    assign data[12061] = 16'b0;
    assign data[12062] = ~16'b0;
    assign data[12063] = ~16'b0;
    assign data[12064] = ~16'b0;
    assign data[12065] = ~16'b0;
    assign data[12066] = ~16'b0;
    assign data[12067] = ~16'b0;
    assign data[12068] = ~16'b0;
    assign data[12069] = ~16'b0;
    assign data[12070] = 16'b0;
    assign data[12071] = 16'b0;
    assign data[12072] = ~16'b0;
    assign data[12073] = ~16'b0;
    assign data[12074] = ~16'b0;
    assign data[12075] = ~16'b0;
    assign data[12076] = ~16'b0;
    assign data[12077] = ~16'b0;
    assign data[12078] = ~16'b0;
    assign data[12079] = ~16'b0;
    assign data[12080] = 16'b0;
    assign data[12081] = 16'b0;
    assign data[12082] = ~16'b0;
    assign data[12083] = ~16'b0;
    assign data[12084] = ~16'b0;
    assign data[12085] = ~16'b0;
    assign data[12086] = ~16'b0;
    assign data[12087] = ~16'b0;
    assign data[12088] = ~16'b0;
    assign data[12089] = ~16'b0;
    assign data[12090] = 16'b0;
    assign data[12091] = 16'b0;
    assign data[12092] = ~16'b0;
    assign data[12093] = ~16'b0;
    assign data[12094] = ~16'b0;
    assign data[12095] = ~16'b0;
    assign data[12096] = ~16'b0;
    assign data[12097] = ~16'b0;
    assign data[12098] = ~16'b0;
    assign data[12099] = ~16'b0;
    assign data[12100] = 16'b0;
    assign data[12101] = 16'b0;
    assign data[12102] = ~16'b0;
    assign data[12103] = ~16'b0;
    assign data[12104] = ~16'b0;
    assign data[12105] = ~16'b0;
    assign data[12106] = ~16'b0;
    assign data[12107] = ~16'b0;
    assign data[12108] = ~16'b0;
    assign data[12109] = ~16'b0;
    assign data[12110] = 16'b0;
    assign data[12111] = 16'b0;
    assign data[12112] = ~16'b0;
    assign data[12113] = ~16'b0;
    assign data[12114] = ~16'b0;
    assign data[12115] = ~16'b0;
    assign data[12116] = ~16'b0;
    assign data[12117] = ~16'b0;
    assign data[12118] = ~16'b0;
    assign data[12119] = ~16'b0;
    assign data[12120] = 16'b0;
    assign data[12121] = 16'b0;
    assign data[12122] = ~16'b0;
    assign data[12123] = ~16'b0;
    assign data[12124] = ~16'b0;
    assign data[12125] = ~16'b0;
    assign data[12126] = ~16'b0;
    assign data[12127] = ~16'b0;
    assign data[12128] = ~16'b0;
    assign data[12129] = ~16'b0;
    assign data[12130] = 16'b0;
    assign data[12131] = 16'b0;
    assign data[12132] = ~16'b0;
    assign data[12133] = ~16'b0;
    assign data[12134] = ~16'b0;
    assign data[12135] = ~16'b0;
    assign data[12136] = ~16'b0;
    assign data[12137] = ~16'b0;
    assign data[12138] = ~16'b0;
    assign data[12139] = ~16'b0;
    assign data[12140] = 16'b0;
    assign data[12141] = 16'b0;
    assign data[12142] = ~16'b0;
    assign data[12143] = ~16'b0;
    assign data[12144] = ~16'b0;
    assign data[12145] = ~16'b0;
    assign data[12146] = ~16'b0;
    assign data[12147] = ~16'b0;
    assign data[12148] = ~16'b0;
    assign data[12149] = ~16'b0;
    assign data[12150] = 16'b0;
    assign data[12151] = 16'b0;
    assign data[12152] = ~16'b0;
    assign data[12153] = ~16'b0;
    assign data[12154] = ~16'b0;
    assign data[12155] = ~16'b0;
    assign data[12156] = ~16'b0;
    assign data[12157] = ~16'b0;
    assign data[12158] = ~16'b0;
    assign data[12159] = ~16'b0;
    assign data[12160] = 16'b0;
    assign data[12161] = 16'b0;
    assign data[12162] = ~16'b0;
    assign data[12163] = ~16'b0;
    assign data[12164] = ~16'b0;
    assign data[12165] = ~16'b0;
    assign data[12166] = ~16'b0;
    assign data[12167] = ~16'b0;
    assign data[12168] = ~16'b0;
    assign data[12169] = ~16'b0;
    assign data[12170] = 16'b0;
    assign data[12171] = 16'b0;
    assign data[12172] = ~16'b0;
    assign data[12173] = ~16'b0;
    assign data[12174] = ~16'b0;
    assign data[12175] = ~16'b0;
    assign data[12176] = ~16'b0;
    assign data[12177] = ~16'b0;
    assign data[12178] = ~16'b0;
    assign data[12179] = ~16'b0;
    assign data[12180] = 16'b0;
    assign data[12181] = 16'b0;
    assign data[12182] = ~16'b0;
    assign data[12183] = ~16'b0;
    assign data[12184] = ~16'b0;
    assign data[12185] = ~16'b0;
    assign data[12186] = ~16'b0;
    assign data[12187] = ~16'b0;
    assign data[12188] = ~16'b0;
    assign data[12189] = ~16'b0;
    assign data[12190] = 16'b0;
    assign data[12191] = 16'b0;
    assign data[12192] = ~16'b0;
    assign data[12193] = ~16'b0;
    assign data[12194] = ~16'b0;
    assign data[12195] = ~16'b0;
    assign data[12196] = ~16'b0;
    assign data[12197] = ~16'b0;
    assign data[12198] = ~16'b0;
    assign data[12199] = ~16'b0;
    assign data[12200] = 16'b0;
    assign data[12201] = 16'b0;
    assign data[12202] = ~16'b0;
    assign data[12203] = ~16'b0;
    assign data[12204] = ~16'b0;
    assign data[12205] = ~16'b0;
    assign data[12206] = ~16'b0;
    assign data[12207] = ~16'b0;
    assign data[12208] = ~16'b0;
    assign data[12209] = ~16'b0;
    assign data[12210] = 16'b0;
    assign data[12211] = 16'b0;
    assign data[12212] = ~16'b0;
    assign data[12213] = ~16'b0;
    assign data[12214] = ~16'b0;
    assign data[12215] = ~16'b0;
    assign data[12216] = ~16'b0;
    assign data[12217] = ~16'b0;
    assign data[12218] = ~16'b0;
    assign data[12219] = ~16'b0;
    assign data[12220] = 16'b0;
    assign data[12221] = 16'b0;
    assign data[12222] = ~16'b0;
    assign data[12223] = ~16'b0;
    assign data[12224] = ~16'b0;
    assign data[12225] = ~16'b0;
    assign data[12226] = ~16'b0;
    assign data[12227] = ~16'b0;
    assign data[12228] = ~16'b0;
    assign data[12229] = ~16'b0;
    assign data[12230] = 16'b0;
    assign data[12231] = 16'b0;
    assign data[12232] = ~16'b0;
    assign data[12233] = ~16'b0;
    assign data[12234] = ~16'b0;
    assign data[12235] = ~16'b0;
    assign data[12236] = ~16'b0;
    assign data[12237] = ~16'b0;
    assign data[12238] = ~16'b0;
    assign data[12239] = ~16'b0;
    assign data[12240] = 16'b0;
    assign data[12241] = 16'b0;
    assign data[12242] = 16'b0;
    assign data[12243] = 16'b0;
    assign data[12244] = 16'b0;
    assign data[12245] = 16'b0;
    assign data[12246] = 16'b0;
    assign data[12247] = 16'b0;
    assign data[12248] = 16'b0;
    assign data[12249] = 16'b0;
    assign data[12250] = 16'b0;
    assign data[12251] = 16'b0;
    assign data[12252] = 16'b0;
    assign data[12253] = 16'b0;
    assign data[12254] = 16'b0;
    assign data[12255] = 16'b0;
    assign data[12256] = 16'b0;
    assign data[12257] = 16'b0;
    assign data[12258] = 16'b0;
    assign data[12259] = 16'b0;
    assign data[12260] = ~16'b0;
    assign data[12261] = ~16'b0;
    assign data[12262] = ~16'b0;
    assign data[12263] = ~16'b0;
    assign data[12264] = ~16'b0;
    assign data[12265] = ~16'b0;
    assign data[12266] = ~16'b0;
    assign data[12267] = ~16'b0;
    assign data[12268] = ~16'b0;
    assign data[12269] = ~16'b0;
    assign data[12270] = ~16'b0;
    assign data[12271] = ~16'b0;
    assign data[12272] = ~16'b0;
    assign data[12273] = ~16'b0;
    assign data[12274] = ~16'b0;
    assign data[12275] = ~16'b0;
    assign data[12276] = ~16'b0;
    assign data[12277] = ~16'b0;
    assign data[12278] = ~16'b0;
    assign data[12279] = ~16'b0;
    assign data[12280] = ~16'b0;
    assign data[12281] = ~16'b0;
    assign data[12282] = ~16'b0;
    assign data[12283] = ~16'b0;
    assign data[12284] = ~16'b0;
    assign data[12285] = ~16'b0;
    assign data[12286] = ~16'b0;
    assign data[12287] = ~16'b0;
    assign data[12288] = ~16'b0;
    assign data[12289] = ~16'b0;
    assign data[12290] = ~16'b0;
    assign data[12291] = ~16'b0;
    assign data[12292] = ~16'b0;
    assign data[12293] = ~16'b0;
    assign data[12294] = ~16'b0;
    assign data[12295] = ~16'b0;
    assign data[12296] = ~16'b0;
    assign data[12297] = ~16'b0;
    assign data[12298] = ~16'b0;
    assign data[12299] = ~16'b0;
    assign data[12300] = ~16'b0;
    assign data[12301] = ~16'b0;
    assign data[12302] = ~16'b0;
    assign data[12303] = ~16'b0;
    assign data[12304] = ~16'b0;
    assign data[12305] = ~16'b0;
    assign data[12306] = ~16'b0;
    assign data[12307] = ~16'b0;
    assign data[12308] = ~16'b0;
    assign data[12309] = ~16'b0;
    assign data[12310] = ~16'b0;
    assign data[12311] = ~16'b0;
    assign data[12312] = ~16'b0;
    assign data[12313] = ~16'b0;
    assign data[12314] = ~16'b0;
    assign data[12315] = ~16'b0;
    assign data[12316] = ~16'b0;
    assign data[12317] = ~16'b0;
    assign data[12318] = ~16'b0;
    assign data[12319] = ~16'b0;
    assign data[12320] = ~16'b0;
    assign data[12321] = ~16'b0;
    assign data[12322] = ~16'b0;
    assign data[12323] = ~16'b0;
    assign data[12324] = ~16'b0;
    assign data[12325] = ~16'b0;
    assign data[12326] = ~16'b0;
    assign data[12327] = ~16'b0;
    assign data[12328] = ~16'b0;
    assign data[12329] = ~16'b0;
    assign data[12330] = ~16'b0;
    assign data[12331] = ~16'b0;
    assign data[12332] = ~16'b0;
    assign data[12333] = ~16'b0;
    assign data[12334] = ~16'b0;
    assign data[12335] = ~16'b0;
    assign data[12336] = ~16'b0;
    assign data[12337] = ~16'b0;
    assign data[12338] = ~16'b0;
    assign data[12339] = ~16'b0;
    assign data[12340] = ~16'b0;
    assign data[12341] = ~16'b0;
    assign data[12342] = ~16'b0;
    assign data[12343] = ~16'b0;
    assign data[12344] = ~16'b0;
    assign data[12345] = ~16'b0;
    assign data[12346] = ~16'b0;
    assign data[12347] = ~16'b0;
    assign data[12348] = ~16'b0;
    assign data[12349] = ~16'b0;
    assign data[12350] = ~16'b0;
    assign data[12351] = ~16'b0;
    assign data[12352] = ~16'b0;
    assign data[12353] = ~16'b0;
    assign data[12354] = ~16'b0;
    assign data[12355] = ~16'b0;
    assign data[12356] = ~16'b0;
    assign data[12357] = ~16'b0;
    assign data[12358] = ~16'b0;
    assign data[12359] = ~16'b0;
    assign data[12360] = ~16'b0;
    assign data[12361] = ~16'b0;
    assign data[12362] = ~16'b0;
    assign data[12363] = ~16'b0;
    assign data[12364] = ~16'b0;
    assign data[12365] = ~16'b0;
    assign data[12366] = ~16'b0;
    assign data[12367] = ~16'b0;
    assign data[12368] = ~16'b0;
    assign data[12369] = ~16'b0;
    assign data[12370] = ~16'b0;
    assign data[12371] = ~16'b0;
    assign data[12372] = ~16'b0;
    assign data[12373] = ~16'b0;
    assign data[12374] = ~16'b0;
    assign data[12375] = ~16'b0;
    assign data[12376] = ~16'b0;
    assign data[12377] = ~16'b0;
    assign data[12378] = ~16'b0;
    assign data[12379] = ~16'b0;
    assign data[12380] = ~16'b0;
    assign data[12381] = ~16'b0;
    assign data[12382] = ~16'b0;
    assign data[12383] = ~16'b0;
    assign data[12384] = ~16'b0;
    assign data[12385] = ~16'b0;
    assign data[12386] = ~16'b0;
    assign data[12387] = ~16'b0;
    assign data[12388] = ~16'b0;
    assign data[12389] = ~16'b0;
    assign data[12390] = ~16'b0;
    assign data[12391] = ~16'b0;
    assign data[12392] = ~16'b0;
    assign data[12393] = ~16'b0;
    assign data[12394] = ~16'b0;
    assign data[12395] = ~16'b0;
    assign data[12396] = ~16'b0;
    assign data[12397] = ~16'b0;
    assign data[12398] = ~16'b0;
    assign data[12399] = ~16'b0;
    assign data[12400] = 16'b0;
    assign data[12401] = 16'b0;
    assign data[12402] = 16'b0;
    assign data[12403] = 16'b0;
    assign data[12404] = 16'b0;
    assign data[12405] = 16'b0;
    assign data[12406] = 16'b0;
    assign data[12407] = 16'b0;
    assign data[12408] = 16'b0;
    assign data[12409] = 16'b0;
    assign data[12410] = 16'b0;
    assign data[12411] = 16'b0;
    assign data[12412] = 16'b0;
    assign data[12413] = 16'b0;
    assign data[12414] = 16'b0;
    assign data[12415] = 16'b0;
    assign data[12416] = 16'b0;
    assign data[12417] = 16'b0;
    assign data[12418] = 16'b0;
    assign data[12419] = 16'b0;
    assign data[12420] = 16'b0;
    assign data[12421] = 16'b0;
    assign data[12422] = ~16'b0;
    assign data[12423] = ~16'b0;
    assign data[12424] = ~16'b0;
    assign data[12425] = ~16'b0;
    assign data[12426] = ~16'b0;
    assign data[12427] = ~16'b0;
    assign data[12428] = ~16'b0;
    assign data[12429] = ~16'b0;
    assign data[12430] = 16'b0;
    assign data[12431] = 16'b0;
    assign data[12432] = ~16'b0;
    assign data[12433] = ~16'b0;
    assign data[12434] = ~16'b0;
    assign data[12435] = ~16'b0;
    assign data[12436] = ~16'b0;
    assign data[12437] = ~16'b0;
    assign data[12438] = ~16'b0;
    assign data[12439] = ~16'b0;
    assign data[12440] = 16'b0;
    assign data[12441] = 16'b0;
    assign data[12442] = ~16'b0;
    assign data[12443] = ~16'b0;
    assign data[12444] = ~16'b0;
    assign data[12445] = ~16'b0;
    assign data[12446] = ~16'b0;
    assign data[12447] = ~16'b0;
    assign data[12448] = ~16'b0;
    assign data[12449] = ~16'b0;
    assign data[12450] = 16'b0;
    assign data[12451] = 16'b0;
    assign data[12452] = ~16'b0;
    assign data[12453] = ~16'b0;
    assign data[12454] = ~16'b0;
    assign data[12455] = ~16'b0;
    assign data[12456] = ~16'b0;
    assign data[12457] = ~16'b0;
    assign data[12458] = ~16'b0;
    assign data[12459] = ~16'b0;
    assign data[12460] = 16'b0;
    assign data[12461] = 16'b0;
    assign data[12462] = ~16'b0;
    assign data[12463] = ~16'b0;
    assign data[12464] = ~16'b0;
    assign data[12465] = ~16'b0;
    assign data[12466] = ~16'b0;
    assign data[12467] = ~16'b0;
    assign data[12468] = ~16'b0;
    assign data[12469] = ~16'b0;
    assign data[12470] = 16'b0;
    assign data[12471] = 16'b0;
    assign data[12472] = ~16'b0;
    assign data[12473] = ~16'b0;
    assign data[12474] = ~16'b0;
    assign data[12475] = ~16'b0;
    assign data[12476] = ~16'b0;
    assign data[12477] = ~16'b0;
    assign data[12478] = ~16'b0;
    assign data[12479] = ~16'b0;
    assign data[12480] = 16'b0;
    assign data[12481] = 16'b0;
    assign data[12482] = ~16'b0;
    assign data[12483] = ~16'b0;
    assign data[12484] = ~16'b0;
    assign data[12485] = ~16'b0;
    assign data[12486] = ~16'b0;
    assign data[12487] = ~16'b0;
    assign data[12488] = ~16'b0;
    assign data[12489] = ~16'b0;
    assign data[12490] = 16'b0;
    assign data[12491] = 16'b0;
    assign data[12492] = ~16'b0;
    assign data[12493] = ~16'b0;
    assign data[12494] = ~16'b0;
    assign data[12495] = ~16'b0;
    assign data[12496] = ~16'b0;
    assign data[12497] = ~16'b0;
    assign data[12498] = ~16'b0;
    assign data[12499] = ~16'b0;
    assign data[12500] = 16'b0;
    assign data[12501] = 16'b0;
    assign data[12502] = ~16'b0;
    assign data[12503] = ~16'b0;
    assign data[12504] = ~16'b0;
    assign data[12505] = ~16'b0;
    assign data[12506] = ~16'b0;
    assign data[12507] = ~16'b0;
    assign data[12508] = ~16'b0;
    assign data[12509] = ~16'b0;
    assign data[12510] = 16'b0;
    assign data[12511] = 16'b0;
    assign data[12512] = ~16'b0;
    assign data[12513] = ~16'b0;
    assign data[12514] = ~16'b0;
    assign data[12515] = ~16'b0;
    assign data[12516] = ~16'b0;
    assign data[12517] = ~16'b0;
    assign data[12518] = ~16'b0;
    assign data[12519] = ~16'b0;
    assign data[12520] = 16'b0;
    assign data[12521] = 16'b0;
    assign data[12522] = ~16'b0;
    assign data[12523] = ~16'b0;
    assign data[12524] = ~16'b0;
    assign data[12525] = ~16'b0;
    assign data[12526] = ~16'b0;
    assign data[12527] = ~16'b0;
    assign data[12528] = ~16'b0;
    assign data[12529] = ~16'b0;
    assign data[12530] = 16'b0;
    assign data[12531] = 16'b0;
    assign data[12532] = ~16'b0;
    assign data[12533] = ~16'b0;
    assign data[12534] = ~16'b0;
    assign data[12535] = ~16'b0;
    assign data[12536] = ~16'b0;
    assign data[12537] = ~16'b0;
    assign data[12538] = ~16'b0;
    assign data[12539] = ~16'b0;
    assign data[12540] = 16'b0;
    assign data[12541] = 16'b0;
    assign data[12542] = ~16'b0;
    assign data[12543] = ~16'b0;
    assign data[12544] = ~16'b0;
    assign data[12545] = ~16'b0;
    assign data[12546] = ~16'b0;
    assign data[12547] = ~16'b0;
    assign data[12548] = ~16'b0;
    assign data[12549] = ~16'b0;
    assign data[12550] = 16'b0;
    assign data[12551] = 16'b0;
    assign data[12552] = ~16'b0;
    assign data[12553] = ~16'b0;
    assign data[12554] = ~16'b0;
    assign data[12555] = ~16'b0;
    assign data[12556] = ~16'b0;
    assign data[12557] = ~16'b0;
    assign data[12558] = ~16'b0;
    assign data[12559] = ~16'b0;
    assign data[12560] = 16'b0;
    assign data[12561] = 16'b0;
    assign data[12562] = ~16'b0;
    assign data[12563] = ~16'b0;
    assign data[12564] = ~16'b0;
    assign data[12565] = ~16'b0;
    assign data[12566] = ~16'b0;
    assign data[12567] = ~16'b0;
    assign data[12568] = ~16'b0;
    assign data[12569] = ~16'b0;
    assign data[12570] = 16'b0;
    assign data[12571] = 16'b0;
    assign data[12572] = ~16'b0;
    assign data[12573] = ~16'b0;
    assign data[12574] = ~16'b0;
    assign data[12575] = ~16'b0;
    assign data[12576] = ~16'b0;
    assign data[12577] = ~16'b0;
    assign data[12578] = ~16'b0;
    assign data[12579] = ~16'b0;
    assign data[12580] = 16'b0;
    assign data[12581] = 16'b0;
    assign data[12582] = ~16'b0;
    assign data[12583] = ~16'b0;
    assign data[12584] = ~16'b0;
    assign data[12585] = ~16'b0;
    assign data[12586] = ~16'b0;
    assign data[12587] = ~16'b0;
    assign data[12588] = ~16'b0;
    assign data[12589] = ~16'b0;
    assign data[12590] = 16'b0;
    assign data[12591] = 16'b0;
    assign data[12592] = ~16'b0;
    assign data[12593] = ~16'b0;
    assign data[12594] = ~16'b0;
    assign data[12595] = ~16'b0;
    assign data[12596] = ~16'b0;
    assign data[12597] = ~16'b0;
    assign data[12598] = ~16'b0;
    assign data[12599] = ~16'b0;
    assign data[12600] = 16'b0;
    assign data[12601] = 16'b0;
    assign data[12602] = ~16'b0;
    assign data[12603] = ~16'b0;
    assign data[12604] = ~16'b0;
    assign data[12605] = ~16'b0;
    assign data[12606] = ~16'b0;
    assign data[12607] = ~16'b0;
    assign data[12608] = ~16'b0;
    assign data[12609] = ~16'b0;
    assign data[12610] = 16'b0;
    assign data[12611] = 16'b0;
    assign data[12612] = ~16'b0;
    assign data[12613] = ~16'b0;
    assign data[12614] = ~16'b0;
    assign data[12615] = ~16'b0;
    assign data[12616] = ~16'b0;
    assign data[12617] = ~16'b0;
    assign data[12618] = ~16'b0;
    assign data[12619] = ~16'b0;
    assign data[12620] = 16'b0;
    assign data[12621] = 16'b0;
    assign data[12622] = ~16'b0;
    assign data[12623] = ~16'b0;
    assign data[12624] = ~16'b0;
    assign data[12625] = ~16'b0;
    assign data[12626] = ~16'b0;
    assign data[12627] = ~16'b0;
    assign data[12628] = ~16'b0;
    assign data[12629] = ~16'b0;
    assign data[12630] = 16'b0;
    assign data[12631] = 16'b0;
    assign data[12632] = ~16'b0;
    assign data[12633] = ~16'b0;
    assign data[12634] = ~16'b0;
    assign data[12635] = ~16'b0;
    assign data[12636] = ~16'b0;
    assign data[12637] = ~16'b0;
    assign data[12638] = ~16'b0;
    assign data[12639] = ~16'b0;
    assign data[12640] = 16'b0;
    assign data[12641] = 16'b0;
    assign data[12642] = ~16'b0;
    assign data[12643] = ~16'b0;
    assign data[12644] = ~16'b0;
    assign data[12645] = ~16'b0;
    assign data[12646] = ~16'b0;
    assign data[12647] = ~16'b0;
    assign data[12648] = ~16'b0;
    assign data[12649] = ~16'b0;
    assign data[12650] = 16'b0;
    assign data[12651] = 16'b0;
    assign data[12652] = ~16'b0;
    assign data[12653] = ~16'b0;
    assign data[12654] = ~16'b0;
    assign data[12655] = ~16'b0;
    assign data[12656] = ~16'b0;
    assign data[12657] = ~16'b0;
    assign data[12658] = ~16'b0;
    assign data[12659] = ~16'b0;
    assign data[12660] = 16'b0;
    assign data[12661] = 16'b0;
    assign data[12662] = ~16'b0;
    assign data[12663] = ~16'b0;
    assign data[12664] = ~16'b0;
    assign data[12665] = ~16'b0;
    assign data[12666] = ~16'b0;
    assign data[12667] = ~16'b0;
    assign data[12668] = ~16'b0;
    assign data[12669] = ~16'b0;
    assign data[12670] = 16'b0;
    assign data[12671] = 16'b0;
    assign data[12672] = ~16'b0;
    assign data[12673] = ~16'b0;
    assign data[12674] = ~16'b0;
    assign data[12675] = ~16'b0;
    assign data[12676] = ~16'b0;
    assign data[12677] = ~16'b0;
    assign data[12678] = ~16'b0;
    assign data[12679] = ~16'b0;
    assign data[12680] = 16'b0;
    assign data[12681] = 16'b0;
    assign data[12682] = ~16'b0;
    assign data[12683] = ~16'b0;
    assign data[12684] = ~16'b0;
    assign data[12685] = ~16'b0;
    assign data[12686] = ~16'b0;
    assign data[12687] = ~16'b0;
    assign data[12688] = ~16'b0;
    assign data[12689] = ~16'b0;
    assign data[12690] = 16'b0;
    assign data[12691] = 16'b0;
    assign data[12692] = ~16'b0;
    assign data[12693] = ~16'b0;
    assign data[12694] = ~16'b0;
    assign data[12695] = ~16'b0;
    assign data[12696] = ~16'b0;
    assign data[12697] = ~16'b0;
    assign data[12698] = ~16'b0;
    assign data[12699] = ~16'b0;
    assign data[12700] = 16'b0;
    assign data[12701] = 16'b0;
    assign data[12702] = ~16'b0;
    assign data[12703] = ~16'b0;
    assign data[12704] = ~16'b0;
    assign data[12705] = ~16'b0;
    assign data[12706] = ~16'b0;
    assign data[12707] = ~16'b0;
    assign data[12708] = ~16'b0;
    assign data[12709] = ~16'b0;
    assign data[12710] = 16'b0;
    assign data[12711] = 16'b0;
    assign data[12712] = ~16'b0;
    assign data[12713] = ~16'b0;
    assign data[12714] = ~16'b0;
    assign data[12715] = ~16'b0;
    assign data[12716] = ~16'b0;
    assign data[12717] = ~16'b0;
    assign data[12718] = ~16'b0;
    assign data[12719] = ~16'b0;
    assign data[12720] = 16'b0;
    assign data[12721] = 16'b0;
    assign data[12722] = ~16'b0;
    assign data[12723] = ~16'b0;
    assign data[12724] = ~16'b0;
    assign data[12725] = ~16'b0;
    assign data[12726] = ~16'b0;
    assign data[12727] = ~16'b0;
    assign data[12728] = ~16'b0;
    assign data[12729] = ~16'b0;
    assign data[12730] = 16'b0;
    assign data[12731] = 16'b0;
    assign data[12732] = ~16'b0;
    assign data[12733] = ~16'b0;
    assign data[12734] = ~16'b0;
    assign data[12735] = ~16'b0;
    assign data[12736] = ~16'b0;
    assign data[12737] = ~16'b0;
    assign data[12738] = ~16'b0;
    assign data[12739] = ~16'b0;
    assign data[12740] = 16'b0;
    assign data[12741] = 16'b0;
    assign data[12742] = ~16'b0;
    assign data[12743] = ~16'b0;
    assign data[12744] = ~16'b0;
    assign data[12745] = ~16'b0;
    assign data[12746] = ~16'b0;
    assign data[12747] = ~16'b0;
    assign data[12748] = ~16'b0;
    assign data[12749] = ~16'b0;
    assign data[12750] = 16'b0;
    assign data[12751] = 16'b0;
    assign data[12752] = ~16'b0;
    assign data[12753] = ~16'b0;
    assign data[12754] = ~16'b0;
    assign data[12755] = ~16'b0;
    assign data[12756] = ~16'b0;
    assign data[12757] = ~16'b0;
    assign data[12758] = ~16'b0;
    assign data[12759] = ~16'b0;
    assign data[12760] = 16'b0;
    assign data[12761] = 16'b0;
    assign data[12762] = ~16'b0;
    assign data[12763] = ~16'b0;
    assign data[12764] = ~16'b0;
    assign data[12765] = ~16'b0;
    assign data[12766] = ~16'b0;
    assign data[12767] = ~16'b0;
    assign data[12768] = ~16'b0;
    assign data[12769] = ~16'b0;
    assign data[12770] = 16'b0;
    assign data[12771] = 16'b0;
    assign data[12772] = 16'b0;
    assign data[12773] = 16'b0;
    assign data[12774] = 16'b0;
    assign data[12775] = 16'b0;
    assign data[12776] = 16'b0;
    assign data[12777] = 16'b0;
    assign data[12778] = 16'b0;
    assign data[12779] = 16'b0;
    assign data[12780] = 16'b0;
    assign data[12781] = 16'b0;
    assign data[12782] = 16'b0;
    assign data[12783] = 16'b0;
    assign data[12784] = 16'b0;
    assign data[12785] = 16'b0;
    assign data[12786] = 16'b0;
    assign data[12787] = 16'b0;
    assign data[12788] = 16'b0;
    assign data[12789] = 16'b0;
    assign data[12790] = ~16'b0;
    assign data[12791] = ~16'b0;
    assign data[12792] = ~16'b0;
    assign data[12793] = ~16'b0;
    assign data[12794] = ~16'b0;
    assign data[12795] = ~16'b0;
    assign data[12796] = ~16'b0;
    assign data[12797] = ~16'b0;
    assign data[12798] = ~16'b0;
    assign data[12799] = ~16'b0;
    assign data[12800] = ~16'b0;
    assign data[12801] = ~16'b0;
    assign data[12802] = ~16'b0;
    assign data[12803] = ~16'b0;
    assign data[12804] = ~16'b0;
    assign data[12805] = ~16'b0;
    assign data[12806] = ~16'b0;
    assign data[12807] = ~16'b0;
    assign data[12808] = ~16'b0;
    assign data[12809] = ~16'b0;
    assign data[12810] = ~16'b0;
    assign data[12811] = ~16'b0;
    assign data[12812] = ~16'b0;
    assign data[12813] = ~16'b0;
    assign data[12814] = ~16'b0;
    assign data[12815] = ~16'b0;
    assign data[12816] = ~16'b0;
    assign data[12817] = ~16'b0;
    assign data[12818] = ~16'b0;
    assign data[12819] = ~16'b0;
    assign data[12820] = ~16'b0;
    assign data[12821] = ~16'b0;
    assign data[12822] = ~16'b0;
    assign data[12823] = ~16'b0;
    assign data[12824] = ~16'b0;
    assign data[12825] = ~16'b0;
    assign data[12826] = ~16'b0;
    assign data[12827] = ~16'b0;
    assign data[12828] = ~16'b0;
    assign data[12829] = ~16'b0;
    assign data[12830] = ~16'b0;
    assign data[12831] = ~16'b0;
    assign data[12832] = ~16'b0;
    assign data[12833] = ~16'b0;
    assign data[12834] = ~16'b0;
    assign data[12835] = ~16'b0;
    assign data[12836] = ~16'b0;
    assign data[12837] = ~16'b0;
    assign data[12838] = ~16'b0;
    assign data[12839] = ~16'b0;
    assign data[12840] = ~16'b0;
    assign data[12841] = ~16'b0;
    assign data[12842] = ~16'b0;
    assign data[12843] = ~16'b0;
    assign data[12844] = ~16'b0;
    assign data[12845] = ~16'b0;
    assign data[12846] = ~16'b0;
    assign data[12847] = ~16'b0;
    assign data[12848] = ~16'b0;
    assign data[12849] = ~16'b0;
    assign data[12850] = ~16'b0;
    assign data[12851] = ~16'b0;
    assign data[12852] = ~16'b0;
    assign data[12853] = ~16'b0;
    assign data[12854] = ~16'b0;
    assign data[12855] = ~16'b0;
    assign data[12856] = ~16'b0;
    assign data[12857] = ~16'b0;
    assign data[12858] = ~16'b0;
    assign data[12859] = ~16'b0;
    assign data[12860] = ~16'b0;
    assign data[12861] = ~16'b0;
    assign data[12862] = ~16'b0;
    assign data[12863] = ~16'b0;
    assign data[12864] = ~16'b0;
    assign data[12865] = ~16'b0;
    assign data[12866] = ~16'b0;
    assign data[12867] = ~16'b0;
    assign data[12868] = ~16'b0;
    assign data[12869] = ~16'b0;
    assign data[12870] = ~16'b0;
    assign data[12871] = ~16'b0;
    assign data[12872] = ~16'b0;
    assign data[12873] = ~16'b0;
    assign data[12874] = ~16'b0;
    assign data[12875] = ~16'b0;
    assign data[12876] = ~16'b0;
    assign data[12877] = ~16'b0;
    assign data[12878] = ~16'b0;
    assign data[12879] = ~16'b0;
    assign data[12880] = ~16'b0;
    assign data[12881] = ~16'b0;
    assign data[12882] = ~16'b0;
    assign data[12883] = ~16'b0;
    assign data[12884] = ~16'b0;
    assign data[12885] = ~16'b0;
    assign data[12886] = ~16'b0;
    assign data[12887] = ~16'b0;
    assign data[12888] = ~16'b0;
    assign data[12889] = ~16'b0;
    assign data[12890] = ~16'b0;
    assign data[12891] = ~16'b0;
    assign data[12892] = ~16'b0;
    assign data[12893] = ~16'b0;
    assign data[12894] = ~16'b0;
    assign data[12895] = ~16'b0;
    assign data[12896] = ~16'b0;
    assign data[12897] = ~16'b0;
    assign data[12898] = ~16'b0;
    assign data[12899] = ~16'b0;
    assign data[12900] = ~16'b0;
    assign data[12901] = ~16'b0;
    assign data[12902] = ~16'b0;
    assign data[12903] = ~16'b0;
    assign data[12904] = ~16'b0;
    assign data[12905] = ~16'b0;
    assign data[12906] = ~16'b0;
    assign data[12907] = ~16'b0;
    assign data[12908] = ~16'b0;
    assign data[12909] = ~16'b0;
    assign data[12910] = ~16'b0;
    assign data[12911] = ~16'b0;
    assign data[12912] = ~16'b0;
    assign data[12913] = ~16'b0;
    assign data[12914] = ~16'b0;
    assign data[12915] = ~16'b0;
    assign data[12916] = ~16'b0;
    assign data[12917] = ~16'b0;
    assign data[12918] = ~16'b0;
    assign data[12919] = ~16'b0;
    assign data[12920] = ~16'b0;
    assign data[12921] = ~16'b0;
    assign data[12922] = ~16'b0;
    assign data[12923] = ~16'b0;
    assign data[12924] = ~16'b0;
    assign data[12925] = ~16'b0;
    assign data[12926] = ~16'b0;
    assign data[12927] = ~16'b0;
    assign data[12928] = ~16'b0;
    assign data[12929] = ~16'b0;
    assign data[12930] = ~16'b0;
    assign data[12931] = ~16'b0;
    assign data[12932] = ~16'b0;
    assign data[12933] = ~16'b0;
    assign data[12934] = ~16'b0;
    assign data[12935] = ~16'b0;
    assign data[12936] = ~16'b0;
    assign data[12937] = ~16'b0;
    assign data[12938] = ~16'b0;
    assign data[12939] = ~16'b0;
    assign data[12940] = ~16'b0;
    assign data[12941] = ~16'b0;
    assign data[12942] = ~16'b0;
    assign data[12943] = ~16'b0;
    assign data[12944] = ~16'b0;
    assign data[12945] = ~16'b0;
    assign data[12946] = ~16'b0;
    assign data[12947] = ~16'b0;
    assign data[12948] = ~16'b0;
    assign data[12949] = ~16'b0;
    assign data[12950] = ~16'b0;
    assign data[12951] = ~16'b0;
    assign data[12952] = ~16'b0;
    assign data[12953] = ~16'b0;
    assign data[12954] = ~16'b0;
    assign data[12955] = ~16'b0;
    assign data[12956] = ~16'b0;
    assign data[12957] = ~16'b0;
    assign data[12958] = ~16'b0;
    assign data[12959] = ~16'b0;
    assign data[12960] = ~16'b0;
    assign data[12961] = ~16'b0;
    assign data[12962] = ~16'b0;
    assign data[12963] = ~16'b0;
    assign data[12964] = ~16'b0;
    assign data[12965] = ~16'b0;
    assign data[12966] = ~16'b0;
    assign data[12967] = ~16'b0;
    assign data[12968] = ~16'b0;
    assign data[12969] = ~16'b0;
    assign data[12970] = ~16'b0;
    assign data[12971] = ~16'b0;
    assign data[12972] = ~16'b0;
    assign data[12973] = ~16'b0;
    assign data[12974] = ~16'b0;
    assign data[12975] = ~16'b0;
    assign data[12976] = ~16'b0;
    assign data[12977] = ~16'b0;
    assign data[12978] = ~16'b0;
    assign data[12979] = ~16'b0;
    assign data[12980] = 16'b0;
    assign data[12981] = 16'b0;
    assign data[12982] = 16'b0;
    assign data[12983] = 16'b0;
    assign data[12984] = 16'b0;
    assign data[12985] = 16'b0;
    assign data[12986] = 16'b0;
    assign data[12987] = 16'b0;
    assign data[12988] = 16'b0;
    assign data[12989] = 16'b0;
    assign data[12990] = 16'b0;
    assign data[12991] = 16'b0;
    assign data[12992] = 16'b0;
    assign data[12993] = 16'b0;
    assign data[12994] = 16'b0;
    assign data[12995] = 16'b0;
    assign data[12996] = 16'b0;
    assign data[12997] = 16'b0;
    assign data[12998] = 16'b0;
    assign data[12999] = 16'b0;
    assign data[13000] = 16'b0;
    assign data[13001] = 16'b0;
    assign data[13002] = ~16'b0;
    assign data[13003] = ~16'b0;
    assign data[13004] = ~16'b0;
    assign data[13005] = ~16'b0;
    assign data[13006] = ~16'b0;
    assign data[13007] = ~16'b0;
    assign data[13008] = ~16'b0;
    assign data[13009] = ~16'b0;
    assign data[13010] = 16'b0;
    assign data[13011] = 16'b0;
    assign data[13012] = ~16'b0;
    assign data[13013] = ~16'b0;
    assign data[13014] = ~16'b0;
    assign data[13015] = ~16'b0;
    assign data[13016] = ~16'b0;
    assign data[13017] = ~16'b0;
    assign data[13018] = ~16'b0;
    assign data[13019] = ~16'b0;
    assign data[13020] = 16'b0;
    assign data[13021] = 16'b0;
    assign data[13022] = ~16'b0;
    assign data[13023] = ~16'b0;
    assign data[13024] = ~16'b0;
    assign data[13025] = ~16'b0;
    assign data[13026] = ~16'b0;
    assign data[13027] = ~16'b0;
    assign data[13028] = ~16'b0;
    assign data[13029] = ~16'b0;
    assign data[13030] = 16'b0;
    assign data[13031] = 16'b0;
    assign data[13032] = ~16'b0;
    assign data[13033] = ~16'b0;
    assign data[13034] = ~16'b0;
    assign data[13035] = ~16'b0;
    assign data[13036] = ~16'b0;
    assign data[13037] = ~16'b0;
    assign data[13038] = ~16'b0;
    assign data[13039] = ~16'b0;
    assign data[13040] = 16'b0;
    assign data[13041] = 16'b0;
    assign data[13042] = ~16'b0;
    assign data[13043] = ~16'b0;
    assign data[13044] = ~16'b0;
    assign data[13045] = ~16'b0;
    assign data[13046] = ~16'b0;
    assign data[13047] = ~16'b0;
    assign data[13048] = ~16'b0;
    assign data[13049] = ~16'b0;
    assign data[13050] = 16'b0;
    assign data[13051] = 16'b0;
    assign data[13052] = ~16'b0;
    assign data[13053] = ~16'b0;
    assign data[13054] = ~16'b0;
    assign data[13055] = ~16'b0;
    assign data[13056] = ~16'b0;
    assign data[13057] = ~16'b0;
    assign data[13058] = ~16'b0;
    assign data[13059] = ~16'b0;
    assign data[13060] = 16'b0;
    assign data[13061] = 16'b0;
    assign data[13062] = ~16'b0;
    assign data[13063] = ~16'b0;
    assign data[13064] = ~16'b0;
    assign data[13065] = ~16'b0;
    assign data[13066] = ~16'b0;
    assign data[13067] = ~16'b0;
    assign data[13068] = ~16'b0;
    assign data[13069] = ~16'b0;
    assign data[13070] = 16'b0;
    assign data[13071] = 16'b0;
    assign data[13072] = ~16'b0;
    assign data[13073] = ~16'b0;
    assign data[13074] = ~16'b0;
    assign data[13075] = ~16'b0;
    assign data[13076] = ~16'b0;
    assign data[13077] = ~16'b0;
    assign data[13078] = ~16'b0;
    assign data[13079] = ~16'b0;
    assign data[13080] = 16'b0;
    assign data[13081] = 16'b0;
    assign data[13082] = ~16'b0;
    assign data[13083] = ~16'b0;
    assign data[13084] = ~16'b0;
    assign data[13085] = ~16'b0;
    assign data[13086] = ~16'b0;
    assign data[13087] = ~16'b0;
    assign data[13088] = ~16'b0;
    assign data[13089] = ~16'b0;
    assign data[13090] = 16'b0;
    assign data[13091] = 16'b0;
    assign data[13092] = ~16'b0;
    assign data[13093] = ~16'b0;
    assign data[13094] = ~16'b0;
    assign data[13095] = ~16'b0;
    assign data[13096] = ~16'b0;
    assign data[13097] = ~16'b0;
    assign data[13098] = ~16'b0;
    assign data[13099] = ~16'b0;
    assign data[13100] = 16'b0;
    assign data[13101] = 16'b0;
    assign data[13102] = ~16'b0;
    assign data[13103] = ~16'b0;
    assign data[13104] = ~16'b0;
    assign data[13105] = ~16'b0;
    assign data[13106] = ~16'b0;
    assign data[13107] = ~16'b0;
    assign data[13108] = ~16'b0;
    assign data[13109] = ~16'b0;
    assign data[13110] = 16'b0;
    assign data[13111] = 16'b0;
    assign data[13112] = ~16'b0;
    assign data[13113] = ~16'b0;
    assign data[13114] = ~16'b0;
    assign data[13115] = ~16'b0;
    assign data[13116] = ~16'b0;
    assign data[13117] = ~16'b0;
    assign data[13118] = ~16'b0;
    assign data[13119] = ~16'b0;
    assign data[13120] = 16'b0;
    assign data[13121] = 16'b0;
    assign data[13122] = ~16'b0;
    assign data[13123] = ~16'b0;
    assign data[13124] = ~16'b0;
    assign data[13125] = ~16'b0;
    assign data[13126] = ~16'b0;
    assign data[13127] = ~16'b0;
    assign data[13128] = ~16'b0;
    assign data[13129] = ~16'b0;
    assign data[13130] = 16'b0;
    assign data[13131] = 16'b0;
    assign data[13132] = ~16'b0;
    assign data[13133] = ~16'b0;
    assign data[13134] = ~16'b0;
    assign data[13135] = ~16'b0;
    assign data[13136] = ~16'b0;
    assign data[13137] = ~16'b0;
    assign data[13138] = ~16'b0;
    assign data[13139] = ~16'b0;
    assign data[13140] = 16'b0;
    assign data[13141] = 16'b0;
    assign data[13142] = ~16'b0;
    assign data[13143] = ~16'b0;
    assign data[13144] = ~16'b0;
    assign data[13145] = ~16'b0;
    assign data[13146] = ~16'b0;
    assign data[13147] = ~16'b0;
    assign data[13148] = ~16'b0;
    assign data[13149] = ~16'b0;
    assign data[13150] = 16'b0;
    assign data[13151] = 16'b0;
    assign data[13152] = ~16'b0;
    assign data[13153] = ~16'b0;
    assign data[13154] = ~16'b0;
    assign data[13155] = ~16'b0;
    assign data[13156] = ~16'b0;
    assign data[13157] = ~16'b0;
    assign data[13158] = ~16'b0;
    assign data[13159] = ~16'b0;
    assign data[13160] = 16'b0;
    assign data[13161] = 16'b0;
    assign data[13162] = ~16'b0;
    assign data[13163] = ~16'b0;
    assign data[13164] = ~16'b0;
    assign data[13165] = ~16'b0;
    assign data[13166] = ~16'b0;
    assign data[13167] = ~16'b0;
    assign data[13168] = ~16'b0;
    assign data[13169] = ~16'b0;
    assign data[13170] = 16'b0;
    assign data[13171] = 16'b0;
    assign data[13172] = ~16'b0;
    assign data[13173] = ~16'b0;
    assign data[13174] = ~16'b0;
    assign data[13175] = ~16'b0;
    assign data[13176] = ~16'b0;
    assign data[13177] = ~16'b0;
    assign data[13178] = ~16'b0;
    assign data[13179] = ~16'b0;
    assign data[13180] = 16'b0;
    assign data[13181] = 16'b0;
    assign data[13182] = ~16'b0;
    assign data[13183] = ~16'b0;
    assign data[13184] = ~16'b0;
    assign data[13185] = ~16'b0;
    assign data[13186] = ~16'b0;
    assign data[13187] = ~16'b0;
    assign data[13188] = ~16'b0;
    assign data[13189] = ~16'b0;
    assign data[13190] = 16'b0;
    assign data[13191] = 16'b0;
    assign data[13192] = ~16'b0;
    assign data[13193] = ~16'b0;
    assign data[13194] = ~16'b0;
    assign data[13195] = ~16'b0;
    assign data[13196] = ~16'b0;
    assign data[13197] = ~16'b0;
    assign data[13198] = ~16'b0;
    assign data[13199] = ~16'b0;
    assign data[13200] = 16'b0;
    assign data[13201] = 16'b0;
    assign data[13202] = ~16'b0;
    assign data[13203] = ~16'b0;
    assign data[13204] = ~16'b0;
    assign data[13205] = ~16'b0;
    assign data[13206] = ~16'b0;
    assign data[13207] = ~16'b0;
    assign data[13208] = ~16'b0;
    assign data[13209] = ~16'b0;
    assign data[13210] = 16'b0;
    assign data[13211] = 16'b0;
    assign data[13212] = ~16'b0;
    assign data[13213] = ~16'b0;
    assign data[13214] = ~16'b0;
    assign data[13215] = ~16'b0;
    assign data[13216] = ~16'b0;
    assign data[13217] = ~16'b0;
    assign data[13218] = ~16'b0;
    assign data[13219] = ~16'b0;
    assign data[13220] = 16'b0;
    assign data[13221] = 16'b0;
    assign data[13222] = ~16'b0;
    assign data[13223] = ~16'b0;
    assign data[13224] = ~16'b0;
    assign data[13225] = ~16'b0;
    assign data[13226] = ~16'b0;
    assign data[13227] = ~16'b0;
    assign data[13228] = ~16'b0;
    assign data[13229] = ~16'b0;
    assign data[13230] = 16'b0;
    assign data[13231] = 16'b0;
    assign data[13232] = ~16'b0;
    assign data[13233] = ~16'b0;
    assign data[13234] = ~16'b0;
    assign data[13235] = ~16'b0;
    assign data[13236] = ~16'b0;
    assign data[13237] = ~16'b0;
    assign data[13238] = ~16'b0;
    assign data[13239] = ~16'b0;
    assign data[13240] = 16'b0;
    assign data[13241] = 16'b0;
    assign data[13242] = ~16'b0;
    assign data[13243] = ~16'b0;
    assign data[13244] = ~16'b0;
    assign data[13245] = ~16'b0;
    assign data[13246] = ~16'b0;
    assign data[13247] = ~16'b0;
    assign data[13248] = ~16'b0;
    assign data[13249] = ~16'b0;
    assign data[13250] = 16'b0;
    assign data[13251] = 16'b0;
    assign data[13252] = ~16'b0;
    assign data[13253] = ~16'b0;
    assign data[13254] = ~16'b0;
    assign data[13255] = ~16'b0;
    assign data[13256] = ~16'b0;
    assign data[13257] = ~16'b0;
    assign data[13258] = ~16'b0;
    assign data[13259] = ~16'b0;
    assign data[13260] = 16'b0;
    assign data[13261] = 16'b0;
    assign data[13262] = ~16'b0;
    assign data[13263] = ~16'b0;
    assign data[13264] = ~16'b0;
    assign data[13265] = ~16'b0;
    assign data[13266] = ~16'b0;
    assign data[13267] = ~16'b0;
    assign data[13268] = ~16'b0;
    assign data[13269] = ~16'b0;
    assign data[13270] = 16'b0;
    assign data[13271] = 16'b0;
    assign data[13272] = ~16'b0;
    assign data[13273] = ~16'b0;
    assign data[13274] = ~16'b0;
    assign data[13275] = ~16'b0;
    assign data[13276] = ~16'b0;
    assign data[13277] = ~16'b0;
    assign data[13278] = ~16'b0;
    assign data[13279] = ~16'b0;
    assign data[13280] = 16'b0;
    assign data[13281] = 16'b0;
    assign data[13282] = 16'b0;
    assign data[13283] = 16'b0;
    assign data[13284] = 16'b0;
    assign data[13285] = 16'b0;
    assign data[13286] = 16'b0;
    assign data[13287] = 16'b0;
    assign data[13288] = 16'b0;
    assign data[13289] = 16'b0;
    assign data[13290] = 16'b0;
    assign data[13291] = 16'b0;
    assign data[13292] = 16'b0;
    assign data[13293] = 16'b0;
    assign data[13294] = 16'b0;
    assign data[13295] = 16'b0;
    assign data[13296] = 16'b0;
    assign data[13297] = 16'b0;
    assign data[13298] = 16'b0;
    assign data[13299] = 16'b0;
    assign data[13300] = ~16'b0;
    assign data[13301] = ~16'b0;
    assign data[13302] = ~16'b0;
    assign data[13303] = ~16'b0;
    assign data[13304] = ~16'b0;
    assign data[13305] = ~16'b0;
    assign data[13306] = ~16'b0;
    assign data[13307] = ~16'b0;
    assign data[13308] = ~16'b0;
    assign data[13309] = ~16'b0;
    assign data[13310] = ~16'b0;
    assign data[13311] = ~16'b0;
    assign data[13312] = ~16'b0;
    assign data[13313] = ~16'b0;
    assign data[13314] = ~16'b0;
    assign data[13315] = ~16'b0;
    assign data[13316] = ~16'b0;
    assign data[13317] = ~16'b0;
    assign data[13318] = ~16'b0;
    assign data[13319] = ~16'b0;
    assign data[13320] = ~16'b0;
    assign data[13321] = ~16'b0;
    assign data[13322] = ~16'b0;
    assign data[13323] = ~16'b0;
    assign data[13324] = ~16'b0;
    assign data[13325] = ~16'b0;
    assign data[13326] = ~16'b0;
    assign data[13327] = ~16'b0;
    assign data[13328] = ~16'b0;
    assign data[13329] = ~16'b0;
    assign data[13330] = ~16'b0;
    assign data[13331] = ~16'b0;
    assign data[13332] = ~16'b0;
    assign data[13333] = ~16'b0;
    assign data[13334] = ~16'b0;
    assign data[13335] = ~16'b0;
    assign data[13336] = ~16'b0;
    assign data[13337] = ~16'b0;
    assign data[13338] = ~16'b0;
    assign data[13339] = ~16'b0;
    assign data[13340] = ~16'b0;
    assign data[13341] = ~16'b0;
    assign data[13342] = ~16'b0;
    assign data[13343] = ~16'b0;
    assign data[13344] = ~16'b0;
    assign data[13345] = ~16'b0;
    assign data[13346] = ~16'b0;
    assign data[13347] = ~16'b0;
    assign data[13348] = ~16'b0;
    assign data[13349] = ~16'b0;
    assign data[13350] = ~16'b0;
    assign data[13351] = ~16'b0;
    assign data[13352] = ~16'b0;
    assign data[13353] = ~16'b0;
    assign data[13354] = ~16'b0;
    assign data[13355] = ~16'b0;
    assign data[13356] = ~16'b0;
    assign data[13357] = ~16'b0;
    assign data[13358] = ~16'b0;
    assign data[13359] = ~16'b0;
    assign data[13360] = ~16'b0;
    assign data[13361] = ~16'b0;
    assign data[13362] = ~16'b0;
    assign data[13363] = ~16'b0;
    assign data[13364] = ~16'b0;
    assign data[13365] = ~16'b0;
    assign data[13366] = ~16'b0;
    assign data[13367] = ~16'b0;
    assign data[13368] = ~16'b0;
    assign data[13369] = ~16'b0;
    assign data[13370] = ~16'b0;
    assign data[13371] = ~16'b0;
    assign data[13372] = ~16'b0;
    assign data[13373] = ~16'b0;
    assign data[13374] = ~16'b0;
    assign data[13375] = ~16'b0;
    assign data[13376] = ~16'b0;
    assign data[13377] = ~16'b0;
    assign data[13378] = ~16'b0;
    assign data[13379] = ~16'b0;
    assign data[13380] = ~16'b0;
    assign data[13381] = ~16'b0;
    assign data[13382] = ~16'b0;
    assign data[13383] = ~16'b0;
    assign data[13384] = ~16'b0;
    assign data[13385] = ~16'b0;
    assign data[13386] = ~16'b0;
    assign data[13387] = ~16'b0;
    assign data[13388] = ~16'b0;
    assign data[13389] = ~16'b0;
    assign data[13390] = ~16'b0;
    assign data[13391] = ~16'b0;
    assign data[13392] = ~16'b0;
    assign data[13393] = ~16'b0;
    assign data[13394] = ~16'b0;
    assign data[13395] = ~16'b0;
    assign data[13396] = ~16'b0;
    assign data[13397] = ~16'b0;
    assign data[13398] = ~16'b0;
    assign data[13399] = ~16'b0;
    assign data[13400] = ~16'b0;
    assign data[13401] = ~16'b0;
    assign data[13402] = ~16'b0;
    assign data[13403] = ~16'b0;
    assign data[13404] = ~16'b0;
    assign data[13405] = ~16'b0;
    assign data[13406] = ~16'b0;
    assign data[13407] = ~16'b0;
    assign data[13408] = ~16'b0;
    assign data[13409] = ~16'b0;
    assign data[13410] = 16'b0;
    assign data[13411] = 16'b0;
    assign data[13412] = 16'b0;
    assign data[13413] = 16'b0;
    assign data[13414] = 16'b0;
    assign data[13415] = 16'b0;
    assign data[13416] = 16'b0;
    assign data[13417] = 16'b0;
    assign data[13418] = 16'b0;
    assign data[13419] = 16'b0;
    assign data[13420] = 16'b0;
    assign data[13421] = 16'b0;
    assign data[13422] = 16'b0;
    assign data[13423] = 16'b0;
    assign data[13424] = 16'b0;
    assign data[13425] = 16'b0;
    assign data[13426] = 16'b0;
    assign data[13427] = 16'b0;
    assign data[13428] = 16'b0;
    assign data[13429] = 16'b0;
    assign data[13430] = 16'b0;
    assign data[13431] = 16'b0;
    assign data[13432] = ~16'b0;
    assign data[13433] = ~16'b0;
    assign data[13434] = ~16'b0;
    assign data[13435] = ~16'b0;
    assign data[13436] = ~16'b0;
    assign data[13437] = ~16'b0;
    assign data[13438] = ~16'b0;
    assign data[13439] = ~16'b0;
    assign data[13440] = 16'b0;
    assign data[13441] = 16'b0;
    assign data[13442] = ~16'b0;
    assign data[13443] = ~16'b0;
    assign data[13444] = ~16'b0;
    assign data[13445] = ~16'b0;
    assign data[13446] = ~16'b0;
    assign data[13447] = ~16'b0;
    assign data[13448] = ~16'b0;
    assign data[13449] = ~16'b0;
    assign data[13450] = 16'b0;
    assign data[13451] = 16'b0;
    assign data[13452] = ~16'b0;
    assign data[13453] = ~16'b0;
    assign data[13454] = ~16'b0;
    assign data[13455] = ~16'b0;
    assign data[13456] = ~16'b0;
    assign data[13457] = ~16'b0;
    assign data[13458] = ~16'b0;
    assign data[13459] = ~16'b0;
    assign data[13460] = 16'b0;
    assign data[13461] = 16'b0;
    assign data[13462] = ~16'b0;
    assign data[13463] = ~16'b0;
    assign data[13464] = ~16'b0;
    assign data[13465] = ~16'b0;
    assign data[13466] = ~16'b0;
    assign data[13467] = ~16'b0;
    assign data[13468] = ~16'b0;
    assign data[13469] = ~16'b0;
    assign data[13470] = 16'b0;
    assign data[13471] = 16'b0;
    assign data[13472] = ~16'b0;
    assign data[13473] = ~16'b0;
    assign data[13474] = ~16'b0;
    assign data[13475] = ~16'b0;
    assign data[13476] = ~16'b0;
    assign data[13477] = ~16'b0;
    assign data[13478] = ~16'b0;
    assign data[13479] = ~16'b0;
    assign data[13480] = 16'b0;
    assign data[13481] = 16'b0;
    assign data[13482] = ~16'b0;
    assign data[13483] = ~16'b0;
    assign data[13484] = ~16'b0;
    assign data[13485] = ~16'b0;
    assign data[13486] = ~16'b0;
    assign data[13487] = ~16'b0;
    assign data[13488] = ~16'b0;
    assign data[13489] = ~16'b0;
    assign data[13490] = 16'b0;
    assign data[13491] = 16'b0;
    assign data[13492] = ~16'b0;
    assign data[13493] = ~16'b0;
    assign data[13494] = ~16'b0;
    assign data[13495] = ~16'b0;
    assign data[13496] = ~16'b0;
    assign data[13497] = ~16'b0;
    assign data[13498] = ~16'b0;
    assign data[13499] = ~16'b0;
    assign data[13500] = 16'b0;
    assign data[13501] = 16'b0;
    assign data[13502] = ~16'b0;
    assign data[13503] = ~16'b0;
    assign data[13504] = ~16'b0;
    assign data[13505] = ~16'b0;
    assign data[13506] = ~16'b0;
    assign data[13507] = ~16'b0;
    assign data[13508] = ~16'b0;
    assign data[13509] = ~16'b0;
    assign data[13510] = 16'b0;
    assign data[13511] = 16'b0;
    assign data[13512] = ~16'b0;
    assign data[13513] = ~16'b0;
    assign data[13514] = ~16'b0;
    assign data[13515] = ~16'b0;
    assign data[13516] = ~16'b0;
    assign data[13517] = ~16'b0;
    assign data[13518] = ~16'b0;
    assign data[13519] = ~16'b0;
    assign data[13520] = 16'b0;
    assign data[13521] = 16'b0;
    assign data[13522] = ~16'b0;
    assign data[13523] = ~16'b0;
    assign data[13524] = ~16'b0;
    assign data[13525] = ~16'b0;
    assign data[13526] = ~16'b0;
    assign data[13527] = ~16'b0;
    assign data[13528] = ~16'b0;
    assign data[13529] = ~16'b0;
    assign data[13530] = 16'b0;
    assign data[13531] = 16'b0;
    assign data[13532] = ~16'b0;
    assign data[13533] = ~16'b0;
    assign data[13534] = ~16'b0;
    assign data[13535] = ~16'b0;
    assign data[13536] = ~16'b0;
    assign data[13537] = ~16'b0;
    assign data[13538] = ~16'b0;
    assign data[13539] = ~16'b0;
    assign data[13540] = 16'b0;
    assign data[13541] = 16'b0;
    assign data[13542] = ~16'b0;
    assign data[13543] = ~16'b0;
    assign data[13544] = ~16'b0;
    assign data[13545] = ~16'b0;
    assign data[13546] = ~16'b0;
    assign data[13547] = ~16'b0;
    assign data[13548] = ~16'b0;
    assign data[13549] = ~16'b0;
    assign data[13550] = 16'b0;
    assign data[13551] = 16'b0;
    assign data[13552] = ~16'b0;
    assign data[13553] = ~16'b0;
    assign data[13554] = ~16'b0;
    assign data[13555] = ~16'b0;
    assign data[13556] = ~16'b0;
    assign data[13557] = ~16'b0;
    assign data[13558] = ~16'b0;
    assign data[13559] = ~16'b0;
    assign data[13560] = 16'b0;
    assign data[13561] = 16'b0;
    assign data[13562] = ~16'b0;
    assign data[13563] = ~16'b0;
    assign data[13564] = ~16'b0;
    assign data[13565] = ~16'b0;
    assign data[13566] = ~16'b0;
    assign data[13567] = ~16'b0;
    assign data[13568] = ~16'b0;
    assign data[13569] = ~16'b0;
    assign data[13570] = 16'b0;
    assign data[13571] = 16'b0;
    assign data[13572] = ~16'b0;
    assign data[13573] = ~16'b0;
    assign data[13574] = ~16'b0;
    assign data[13575] = ~16'b0;
    assign data[13576] = ~16'b0;
    assign data[13577] = ~16'b0;
    assign data[13578] = ~16'b0;
    assign data[13579] = ~16'b0;
    assign data[13580] = 16'b0;
    assign data[13581] = 16'b0;
    assign data[13582] = ~16'b0;
    assign data[13583] = ~16'b0;
    assign data[13584] = ~16'b0;
    assign data[13585] = ~16'b0;
    assign data[13586] = ~16'b0;
    assign data[13587] = ~16'b0;
    assign data[13588] = ~16'b0;
    assign data[13589] = ~16'b0;
    assign data[13590] = 16'b0;
    assign data[13591] = 16'b0;
    assign data[13592] = ~16'b0;
    assign data[13593] = ~16'b0;
    assign data[13594] = ~16'b0;
    assign data[13595] = ~16'b0;
    assign data[13596] = ~16'b0;
    assign data[13597] = ~16'b0;
    assign data[13598] = ~16'b0;
    assign data[13599] = ~16'b0;
    assign data[13600] = 16'b0;
    assign data[13601] = 16'b0;
    assign data[13602] = ~16'b0;
    assign data[13603] = ~16'b0;
    assign data[13604] = ~16'b0;
    assign data[13605] = ~16'b0;
    assign data[13606] = ~16'b0;
    assign data[13607] = ~16'b0;
    assign data[13608] = ~16'b0;
    assign data[13609] = ~16'b0;
    assign data[13610] = 16'b0;
    assign data[13611] = 16'b0;
    assign data[13612] = ~16'b0;
    assign data[13613] = ~16'b0;
    assign data[13614] = ~16'b0;
    assign data[13615] = ~16'b0;
    assign data[13616] = ~16'b0;
    assign data[13617] = ~16'b0;
    assign data[13618] = ~16'b0;
    assign data[13619] = ~16'b0;
    assign data[13620] = 16'b0;
    assign data[13621] = 16'b0;
    assign data[13622] = ~16'b0;
    assign data[13623] = ~16'b0;
    assign data[13624] = ~16'b0;
    assign data[13625] = ~16'b0;
    assign data[13626] = ~16'b0;
    assign data[13627] = ~16'b0;
    assign data[13628] = ~16'b0;
    assign data[13629] = ~16'b0;
    assign data[13630] = 16'b0;
    assign data[13631] = 16'b0;
    assign data[13632] = ~16'b0;
    assign data[13633] = ~16'b0;
    assign data[13634] = ~16'b0;
    assign data[13635] = ~16'b0;
    assign data[13636] = ~16'b0;
    assign data[13637] = ~16'b0;
    assign data[13638] = ~16'b0;
    assign data[13639] = ~16'b0;
    assign data[13640] = 16'b0;
    assign data[13641] = 16'b0;
    assign data[13642] = ~16'b0;
    assign data[13643] = ~16'b0;
    assign data[13644] = ~16'b0;
    assign data[13645] = ~16'b0;
    assign data[13646] = ~16'b0;
    assign data[13647] = ~16'b0;
    assign data[13648] = ~16'b0;
    assign data[13649] = ~16'b0;
    assign data[13650] = 16'b0;
    assign data[13651] = 16'b0;
    assign data[13652] = ~16'b0;
    assign data[13653] = ~16'b0;
    assign data[13654] = ~16'b0;
    assign data[13655] = ~16'b0;
    assign data[13656] = ~16'b0;
    assign data[13657] = ~16'b0;
    assign data[13658] = ~16'b0;
    assign data[13659] = ~16'b0;
    assign data[13660] = 16'b0;
    assign data[13661] = 16'b0;
    assign data[13662] = ~16'b0;
    assign data[13663] = ~16'b0;
    assign data[13664] = ~16'b0;
    assign data[13665] = ~16'b0;
    assign data[13666] = ~16'b0;
    assign data[13667] = ~16'b0;
    assign data[13668] = ~16'b0;
    assign data[13669] = ~16'b0;
    assign data[13670] = 16'b0;
    assign data[13671] = 16'b0;
    assign data[13672] = ~16'b0;
    assign data[13673] = ~16'b0;
    assign data[13674] = ~16'b0;
    assign data[13675] = ~16'b0;
    assign data[13676] = ~16'b0;
    assign data[13677] = ~16'b0;
    assign data[13678] = ~16'b0;
    assign data[13679] = ~16'b0;
    assign data[13680] = 16'b0;
    assign data[13681] = 16'b0;
    assign data[13682] = ~16'b0;
    assign data[13683] = ~16'b0;
    assign data[13684] = ~16'b0;
    assign data[13685] = ~16'b0;
    assign data[13686] = ~16'b0;
    assign data[13687] = ~16'b0;
    assign data[13688] = ~16'b0;
    assign data[13689] = ~16'b0;
    assign data[13690] = 16'b0;
    assign data[13691] = 16'b0;
    assign data[13692] = ~16'b0;
    assign data[13693] = ~16'b0;
    assign data[13694] = ~16'b0;
    assign data[13695] = ~16'b0;
    assign data[13696] = ~16'b0;
    assign data[13697] = ~16'b0;
    assign data[13698] = ~16'b0;
    assign data[13699] = ~16'b0;
    assign data[13700] = 16'b0;
    assign data[13701] = 16'b0;
    assign data[13702] = ~16'b0;
    assign data[13703] = ~16'b0;
    assign data[13704] = ~16'b0;
    assign data[13705] = ~16'b0;
    assign data[13706] = ~16'b0;
    assign data[13707] = ~16'b0;
    assign data[13708] = ~16'b0;
    assign data[13709] = ~16'b0;
    assign data[13710] = 16'b0;
    assign data[13711] = 16'b0;
    assign data[13712] = ~16'b0;
    assign data[13713] = ~16'b0;
    assign data[13714] = ~16'b0;
    assign data[13715] = ~16'b0;
    assign data[13716] = ~16'b0;
    assign data[13717] = ~16'b0;
    assign data[13718] = ~16'b0;
    assign data[13719] = ~16'b0;
    assign data[13720] = 16'b0;
    assign data[13721] = 16'b0;
    assign data[13722] = ~16'b0;
    assign data[13723] = ~16'b0;
    assign data[13724] = ~16'b0;
    assign data[13725] = ~16'b0;
    assign data[13726] = ~16'b0;
    assign data[13727] = ~16'b0;
    assign data[13728] = ~16'b0;
    assign data[13729] = ~16'b0;
    assign data[13730] = 16'b0;
    assign data[13731] = 16'b0;
    assign data[13732] = ~16'b0;
    assign data[13733] = ~16'b0;
    assign data[13734] = ~16'b0;
    assign data[13735] = ~16'b0;
    assign data[13736] = ~16'b0;
    assign data[13737] = ~16'b0;
    assign data[13738] = ~16'b0;
    assign data[13739] = ~16'b0;
    assign data[13740] = 16'b0;
    assign data[13741] = 16'b0;
    assign data[13742] = ~16'b0;
    assign data[13743] = ~16'b0;
    assign data[13744] = ~16'b0;
    assign data[13745] = ~16'b0;
    assign data[13746] = ~16'b0;
    assign data[13747] = ~16'b0;
    assign data[13748] = ~16'b0;
    assign data[13749] = ~16'b0;
    assign data[13750] = 16'b0;
    assign data[13751] = 16'b0;
    assign data[13752] = ~16'b0;
    assign data[13753] = ~16'b0;
    assign data[13754] = ~16'b0;
    assign data[13755] = ~16'b0;
    assign data[13756] = ~16'b0;
    assign data[13757] = ~16'b0;
    assign data[13758] = ~16'b0;
    assign data[13759] = ~16'b0;
    assign data[13760] = 16'b0;
    assign data[13761] = 16'b0;
    assign data[13762] = ~16'b0;
    assign data[13763] = ~16'b0;
    assign data[13764] = ~16'b0;
    assign data[13765] = ~16'b0;
    assign data[13766] = ~16'b0;
    assign data[13767] = ~16'b0;
    assign data[13768] = ~16'b0;
    assign data[13769] = ~16'b0;
    assign data[13770] = 16'b0;
    assign data[13771] = 16'b0;
    assign data[13772] = ~16'b0;
    assign data[13773] = ~16'b0;
    assign data[13774] = ~16'b0;
    assign data[13775] = ~16'b0;
    assign data[13776] = ~16'b0;
    assign data[13777] = ~16'b0;
    assign data[13778] = ~16'b0;
    assign data[13779] = ~16'b0;
    assign data[13780] = 16'b0;
    assign data[13781] = 16'b0;
    assign data[13782] = 16'b0;
    assign data[13783] = 16'b0;
    assign data[13784] = 16'b0;
    assign data[13785] = 16'b0;
    assign data[13786] = 16'b0;
    assign data[13787] = 16'b0;
    assign data[13788] = 16'b0;
    assign data[13789] = 16'b0;
    assign data[13790] = 16'b0;
    assign data[13791] = 16'b0;
    assign data[13792] = 16'b0;
    assign data[13793] = 16'b0;
    assign data[13794] = 16'b0;
    assign data[13795] = 16'b0;
    assign data[13796] = 16'b0;
    assign data[13797] = 16'b0;
    assign data[13798] = 16'b0;
    assign data[13799] = 16'b0;
    assign data[13800] = ~16'b0;
    assign data[13801] = ~16'b0;
    assign data[13802] = ~16'b0;
    assign data[13803] = ~16'b0;
    assign data[13804] = ~16'b0;
    assign data[13805] = ~16'b0;
    assign data[13806] = ~16'b0;
    assign data[13807] = ~16'b0;
    assign data[13808] = ~16'b0;
    assign data[13809] = ~16'b0;
    assign data[13810] = ~16'b0;
    assign data[13811] = ~16'b0;
    assign data[13812] = ~16'b0;
    assign data[13813] = ~16'b0;
    assign data[13814] = ~16'b0;
    assign data[13815] = ~16'b0;
    assign data[13816] = ~16'b0;
    assign data[13817] = ~16'b0;
    assign data[13818] = ~16'b0;
    assign data[13819] = ~16'b0;
    assign data[13820] = ~16'b0;
    assign data[13821] = ~16'b0;
    assign data[13822] = ~16'b0;
    assign data[13823] = ~16'b0;
    assign data[13824] = ~16'b0;
    assign data[13825] = ~16'b0;
    assign data[13826] = ~16'b0;
    assign data[13827] = ~16'b0;
    assign data[13828] = ~16'b0;
    assign data[13829] = ~16'b0;
    assign data[13830] = ~16'b0;
    assign data[13831] = ~16'b0;
    assign data[13832] = ~16'b0;
    assign data[13833] = ~16'b0;
    assign data[13834] = ~16'b0;
    assign data[13835] = ~16'b0;
    assign data[13836] = ~16'b0;
    assign data[13837] = ~16'b0;
    assign data[13838] = ~16'b0;
    assign data[13839] = ~16'b0;
    assign data[13840] = ~16'b0;
    assign data[13841] = ~16'b0;
    assign data[13842] = ~16'b0;
    assign data[13843] = ~16'b0;
    assign data[13844] = ~16'b0;
    assign data[13845] = ~16'b0;
    assign data[13846] = ~16'b0;
    assign data[13847] = ~16'b0;
    assign data[13848] = ~16'b0;
    assign data[13849] = ~16'b0;
    assign data[13850] = ~16'b0;
    assign data[13851] = ~16'b0;
    assign data[13852] = ~16'b0;
    assign data[13853] = ~16'b0;
    assign data[13854] = ~16'b0;
    assign data[13855] = ~16'b0;
    assign data[13856] = ~16'b0;
    assign data[13857] = ~16'b0;
    assign data[13858] = ~16'b0;
    assign data[13859] = ~16'b0;
    assign data[13860] = ~16'b0;
    assign data[13861] = ~16'b0;
    assign data[13862] = ~16'b0;
    assign data[13863] = ~16'b0;
    assign data[13864] = ~16'b0;
    assign data[13865] = ~16'b0;
    assign data[13866] = ~16'b0;
    assign data[13867] = ~16'b0;
    assign data[13868] = ~16'b0;
    assign data[13869] = ~16'b0;
    assign data[13870] = ~16'b0;
    assign data[13871] = ~16'b0;
    assign data[13872] = ~16'b0;
    assign data[13873] = ~16'b0;
    assign data[13874] = ~16'b0;
    assign data[13875] = ~16'b0;
    assign data[13876] = ~16'b0;
    assign data[13877] = ~16'b0;
    assign data[13878] = ~16'b0;
    assign data[13879] = ~16'b0;
    assign data[13880] = ~16'b0;
    assign data[13881] = ~16'b0;
    assign data[13882] = ~16'b0;
    assign data[13883] = ~16'b0;
    assign data[13884] = ~16'b0;
    assign data[13885] = ~16'b0;
    assign data[13886] = ~16'b0;
    assign data[13887] = ~16'b0;
    assign data[13888] = ~16'b0;
    assign data[13889] = ~16'b0;
    assign data[13890] = ~16'b0;
    assign data[13891] = ~16'b0;
    assign data[13892] = ~16'b0;
    assign data[13893] = ~16'b0;
    assign data[13894] = ~16'b0;
    assign data[13895] = ~16'b0;
    assign data[13896] = ~16'b0;
    assign data[13897] = ~16'b0;
    assign data[13898] = ~16'b0;
    assign data[13899] = ~16'b0;
    assign data[13900] = 16'b0;
    assign data[13901] = 16'b0;
    assign data[13902] = 16'b0;
    assign data[13903] = 16'b0;
    assign data[13904] = 16'b0;
    assign data[13905] = 16'b0;
    assign data[13906] = 16'b0;
    assign data[13907] = 16'b0;
    assign data[13908] = 16'b0;
    assign data[13909] = 16'b0;
    assign data[13910] = 16'b0;
    assign data[13911] = 16'b0;
    assign data[13912] = 16'b0;
    assign data[13913] = 16'b0;
    assign data[13914] = 16'b0;
    assign data[13915] = 16'b0;
    assign data[13916] = 16'b0;
    assign data[13917] = 16'b0;
    assign data[13918] = 16'b0;
    assign data[13919] = 16'b0;
    assign data[13920] = 16'b0;
    assign data[13921] = 16'b0;
    assign data[13922] = ~16'b0;
    assign data[13923] = ~16'b0;
    assign data[13924] = ~16'b0;
    assign data[13925] = ~16'b0;
    assign data[13926] = ~16'b0;
    assign data[13927] = ~16'b0;
    assign data[13928] = ~16'b0;
    assign data[13929] = ~16'b0;
    assign data[13930] = 16'b0;
    assign data[13931] = 16'b0;
    assign data[13932] = ~16'b0;
    assign data[13933] = ~16'b0;
    assign data[13934] = ~16'b0;
    assign data[13935] = ~16'b0;
    assign data[13936] = ~16'b0;
    assign data[13937] = ~16'b0;
    assign data[13938] = ~16'b0;
    assign data[13939] = ~16'b0;
    assign data[13940] = 16'b0;
    assign data[13941] = 16'b0;
    assign data[13942] = ~16'b0;
    assign data[13943] = ~16'b0;
    assign data[13944] = ~16'b0;
    assign data[13945] = ~16'b0;
    assign data[13946] = ~16'b0;
    assign data[13947] = ~16'b0;
    assign data[13948] = ~16'b0;
    assign data[13949] = ~16'b0;
    assign data[13950] = 16'b0;
    assign data[13951] = 16'b0;
    assign data[13952] = ~16'b0;
    assign data[13953] = ~16'b0;
    assign data[13954] = ~16'b0;
    assign data[13955] = ~16'b0;
    assign data[13956] = ~16'b0;
    assign data[13957] = ~16'b0;
    assign data[13958] = ~16'b0;
    assign data[13959] = ~16'b0;
    assign data[13960] = 16'b0;
    assign data[13961] = 16'b0;
    assign data[13962] = ~16'b0;
    assign data[13963] = ~16'b0;
    assign data[13964] = ~16'b0;
    assign data[13965] = ~16'b0;
    assign data[13966] = ~16'b0;
    assign data[13967] = ~16'b0;
    assign data[13968] = ~16'b0;
    assign data[13969] = ~16'b0;
    assign data[13970] = 16'b0;
    assign data[13971] = 16'b0;
    assign data[13972] = ~16'b0;
    assign data[13973] = ~16'b0;
    assign data[13974] = ~16'b0;
    assign data[13975] = ~16'b0;
    assign data[13976] = ~16'b0;
    assign data[13977] = ~16'b0;
    assign data[13978] = ~16'b0;
    assign data[13979] = ~16'b0;
    assign data[13980] = 16'b0;
    assign data[13981] = 16'b0;
    assign data[13982] = ~16'b0;
    assign data[13983] = ~16'b0;
    assign data[13984] = ~16'b0;
    assign data[13985] = ~16'b0;
    assign data[13986] = ~16'b0;
    assign data[13987] = ~16'b0;
    assign data[13988] = ~16'b0;
    assign data[13989] = ~16'b0;
    assign data[13990] = 16'b0;
    assign data[13991] = 16'b0;
    assign data[13992] = ~16'b0;
    assign data[13993] = ~16'b0;
    assign data[13994] = ~16'b0;
    assign data[13995] = ~16'b0;
    assign data[13996] = ~16'b0;
    assign data[13997] = ~16'b0;
    assign data[13998] = ~16'b0;
    assign data[13999] = ~16'b0;
    assign data[14000] = 16'b0;
    assign data[14001] = 16'b0;
    assign data[14002] = ~16'b0;
    assign data[14003] = ~16'b0;
    assign data[14004] = ~16'b0;
    assign data[14005] = ~16'b0;
    assign data[14006] = ~16'b0;
    assign data[14007] = ~16'b0;
    assign data[14008] = ~16'b0;
    assign data[14009] = ~16'b0;
    assign data[14010] = 16'b0;
    assign data[14011] = 16'b0;
    assign data[14012] = ~16'b0;
    assign data[14013] = ~16'b0;
    assign data[14014] = ~16'b0;
    assign data[14015] = ~16'b0;
    assign data[14016] = ~16'b0;
    assign data[14017] = ~16'b0;
    assign data[14018] = ~16'b0;
    assign data[14019] = ~16'b0;
    assign data[14020] = 16'b0;
    assign data[14021] = 16'b0;
    assign data[14022] = ~16'b0;
    assign data[14023] = ~16'b0;
    assign data[14024] = ~16'b0;
    assign data[14025] = ~16'b0;
    assign data[14026] = ~16'b0;
    assign data[14027] = ~16'b0;
    assign data[14028] = ~16'b0;
    assign data[14029] = ~16'b0;
    assign data[14030] = 16'b0;
    assign data[14031] = 16'b0;
    assign data[14032] = ~16'b0;
    assign data[14033] = ~16'b0;
    assign data[14034] = ~16'b0;
    assign data[14035] = ~16'b0;
    assign data[14036] = ~16'b0;
    assign data[14037] = ~16'b0;
    assign data[14038] = ~16'b0;
    assign data[14039] = ~16'b0;
    assign data[14040] = 16'b0;
    assign data[14041] = 16'b0;
    assign data[14042] = ~16'b0;
    assign data[14043] = ~16'b0;
    assign data[14044] = ~16'b0;
    assign data[14045] = ~16'b0;
    assign data[14046] = ~16'b0;
    assign data[14047] = ~16'b0;
    assign data[14048] = ~16'b0;
    assign data[14049] = ~16'b0;
    assign data[14050] = 16'b0;
    assign data[14051] = 16'b0;
    assign data[14052] = ~16'b0;
    assign data[14053] = ~16'b0;
    assign data[14054] = ~16'b0;
    assign data[14055] = ~16'b0;
    assign data[14056] = ~16'b0;
    assign data[14057] = ~16'b0;
    assign data[14058] = ~16'b0;
    assign data[14059] = ~16'b0;
    assign data[14060] = 16'b0;
    assign data[14061] = 16'b0;
    assign data[14062] = ~16'b0;
    assign data[14063] = ~16'b0;
    assign data[14064] = ~16'b0;
    assign data[14065] = ~16'b0;
    assign data[14066] = ~16'b0;
    assign data[14067] = ~16'b0;
    assign data[14068] = ~16'b0;
    assign data[14069] = ~16'b0;
    assign data[14070] = 16'b0;
    assign data[14071] = 16'b0;
    assign data[14072] = ~16'b0;
    assign data[14073] = ~16'b0;
    assign data[14074] = ~16'b0;
    assign data[14075] = ~16'b0;
    assign data[14076] = ~16'b0;
    assign data[14077] = ~16'b0;
    assign data[14078] = ~16'b0;
    assign data[14079] = ~16'b0;
    assign data[14080] = 16'b0;
    assign data[14081] = 16'b0;
    assign data[14082] = ~16'b0;
    assign data[14083] = ~16'b0;
    assign data[14084] = ~16'b0;
    assign data[14085] = ~16'b0;
    assign data[14086] = ~16'b0;
    assign data[14087] = ~16'b0;
    assign data[14088] = ~16'b0;
    assign data[14089] = ~16'b0;
    assign data[14090] = 16'b0;
    assign data[14091] = 16'b0;
    assign data[14092] = ~16'b0;
    assign data[14093] = ~16'b0;
    assign data[14094] = ~16'b0;
    assign data[14095] = ~16'b0;
    assign data[14096] = ~16'b0;
    assign data[14097] = ~16'b0;
    assign data[14098] = ~16'b0;
    assign data[14099] = ~16'b0;
    assign data[14100] = 16'b0;
    assign data[14101] = 16'b0;
    assign data[14102] = ~16'b0;
    assign data[14103] = ~16'b0;
    assign data[14104] = ~16'b0;
    assign data[14105] = ~16'b0;
    assign data[14106] = ~16'b0;
    assign data[14107] = ~16'b0;
    assign data[14108] = ~16'b0;
    assign data[14109] = ~16'b0;
    assign data[14110] = 16'b0;
    assign data[14111] = 16'b0;
    assign data[14112] = ~16'b0;
    assign data[14113] = ~16'b0;
    assign data[14114] = ~16'b0;
    assign data[14115] = ~16'b0;
    assign data[14116] = ~16'b0;
    assign data[14117] = ~16'b0;
    assign data[14118] = ~16'b0;
    assign data[14119] = ~16'b0;
    assign data[14120] = 16'b0;
    assign data[14121] = 16'b0;
    assign data[14122] = ~16'b0;
    assign data[14123] = ~16'b0;
    assign data[14124] = ~16'b0;
    assign data[14125] = ~16'b0;
    assign data[14126] = ~16'b0;
    assign data[14127] = ~16'b0;
    assign data[14128] = ~16'b0;
    assign data[14129] = ~16'b0;
    assign data[14130] = 16'b0;
    assign data[14131] = 16'b0;
    assign data[14132] = ~16'b0;
    assign data[14133] = ~16'b0;
    assign data[14134] = ~16'b0;
    assign data[14135] = ~16'b0;
    assign data[14136] = ~16'b0;
    assign data[14137] = ~16'b0;
    assign data[14138] = ~16'b0;
    assign data[14139] = ~16'b0;
    assign data[14140] = 16'b0;
    assign data[14141] = 16'b0;
    assign data[14142] = ~16'b0;
    assign data[14143] = ~16'b0;
    assign data[14144] = ~16'b0;
    assign data[14145] = ~16'b0;
    assign data[14146] = ~16'b0;
    assign data[14147] = ~16'b0;
    assign data[14148] = ~16'b0;
    assign data[14149] = ~16'b0;
    assign data[14150] = 16'b0;
    assign data[14151] = 16'b0;
    assign data[14152] = ~16'b0;
    assign data[14153] = ~16'b0;
    assign data[14154] = ~16'b0;
    assign data[14155] = ~16'b0;
    assign data[14156] = ~16'b0;
    assign data[14157] = ~16'b0;
    assign data[14158] = ~16'b0;
    assign data[14159] = ~16'b0;
    assign data[14160] = 16'b0;
    assign data[14161] = 16'b0;
    assign data[14162] = ~16'b0;
    assign data[14163] = ~16'b0;
    assign data[14164] = ~16'b0;
    assign data[14165] = ~16'b0;
    assign data[14166] = ~16'b0;
    assign data[14167] = ~16'b0;
    assign data[14168] = ~16'b0;
    assign data[14169] = ~16'b0;
    assign data[14170] = 16'b0;
    assign data[14171] = 16'b0;
    assign data[14172] = ~16'b0;
    assign data[14173] = ~16'b0;
    assign data[14174] = ~16'b0;
    assign data[14175] = ~16'b0;
    assign data[14176] = ~16'b0;
    assign data[14177] = ~16'b0;
    assign data[14178] = ~16'b0;
    assign data[14179] = ~16'b0;
    assign data[14180] = 16'b0;
    assign data[14181] = 16'b0;
    assign data[14182] = ~16'b0;
    assign data[14183] = ~16'b0;
    assign data[14184] = ~16'b0;
    assign data[14185] = ~16'b0;
    assign data[14186] = ~16'b0;
    assign data[14187] = ~16'b0;
    assign data[14188] = ~16'b0;
    assign data[14189] = ~16'b0;
    assign data[14190] = 16'b0;
    assign data[14191] = 16'b0;
    assign data[14192] = ~16'b0;
    assign data[14193] = ~16'b0;
    assign data[14194] = ~16'b0;
    assign data[14195] = ~16'b0;
    assign data[14196] = ~16'b0;
    assign data[14197] = ~16'b0;
    assign data[14198] = ~16'b0;
    assign data[14199] = ~16'b0;
    assign data[14200] = 16'b0;
    assign data[14201] = 16'b0;
    assign data[14202] = ~16'b0;
    assign data[14203] = ~16'b0;
    assign data[14204] = ~16'b0;
    assign data[14205] = ~16'b0;
    assign data[14206] = ~16'b0;
    assign data[14207] = ~16'b0;
    assign data[14208] = ~16'b0;
    assign data[14209] = ~16'b0;
    assign data[14210] = 16'b0;
    assign data[14211] = 16'b0;
    assign data[14212] = ~16'b0;
    assign data[14213] = ~16'b0;
    assign data[14214] = ~16'b0;
    assign data[14215] = ~16'b0;
    assign data[14216] = ~16'b0;
    assign data[14217] = ~16'b0;
    assign data[14218] = ~16'b0;
    assign data[14219] = ~16'b0;
    assign data[14220] = 16'b0;
    assign data[14221] = 16'b0;
    assign data[14222] = ~16'b0;
    assign data[14223] = ~16'b0;
    assign data[14224] = ~16'b0;
    assign data[14225] = ~16'b0;
    assign data[14226] = ~16'b0;
    assign data[14227] = ~16'b0;
    assign data[14228] = ~16'b0;
    assign data[14229] = ~16'b0;
    assign data[14230] = 16'b0;
    assign data[14231] = 16'b0;
    assign data[14232] = ~16'b0;
    assign data[14233] = ~16'b0;
    assign data[14234] = ~16'b0;
    assign data[14235] = ~16'b0;
    assign data[14236] = ~16'b0;
    assign data[14237] = ~16'b0;
    assign data[14238] = ~16'b0;
    assign data[14239] = ~16'b0;
    assign data[14240] = 16'b0;
    assign data[14241] = 16'b0;
    assign data[14242] = ~16'b0;
    assign data[14243] = ~16'b0;
    assign data[14244] = ~16'b0;
    assign data[14245] = ~16'b0;
    assign data[14246] = ~16'b0;
    assign data[14247] = ~16'b0;
    assign data[14248] = ~16'b0;
    assign data[14249] = ~16'b0;
    assign data[14250] = 16'b0;
    assign data[14251] = 16'b0;
    assign data[14252] = ~16'b0;
    assign data[14253] = ~16'b0;
    assign data[14254] = ~16'b0;
    assign data[14255] = ~16'b0;
    assign data[14256] = ~16'b0;
    assign data[14257] = ~16'b0;
    assign data[14258] = ~16'b0;
    assign data[14259] = ~16'b0;
    assign data[14260] = 16'b0;
    assign data[14261] = 16'b0;
    assign data[14262] = ~16'b0;
    assign data[14263] = ~16'b0;
    assign data[14264] = ~16'b0;
    assign data[14265] = ~16'b0;
    assign data[14266] = ~16'b0;
    assign data[14267] = ~16'b0;
    assign data[14268] = ~16'b0;
    assign data[14269] = ~16'b0;
    assign data[14270] = 16'b0;
    assign data[14271] = 16'b0;
    assign data[14272] = 16'b0;
    assign data[14273] = 16'b0;
    assign data[14274] = 16'b0;
    assign data[14275] = 16'b0;
    assign data[14276] = 16'b0;
    assign data[14277] = 16'b0;
    assign data[14278] = 16'b0;
    assign data[14279] = 16'b0;
    assign data[14280] = 16'b0;
    assign data[14281] = 16'b0;
    assign data[14282] = 16'b0;
    assign data[14283] = 16'b0;
    assign data[14284] = 16'b0;
    assign data[14285] = 16'b0;
    assign data[14286] = 16'b0;
    assign data[14287] = 16'b0;
    assign data[14288] = 16'b0;
    assign data[14289] = 16'b0;
    assign data[14290] = ~16'b0;
    assign data[14291] = ~16'b0;
    assign data[14292] = ~16'b0;
    assign data[14293] = ~16'b0;
    assign data[14294] = ~16'b0;
    assign data[14295] = ~16'b0;
    assign data[14296] = ~16'b0;
    assign data[14297] = ~16'b0;
    assign data[14298] = ~16'b0;
    assign data[14299] = ~16'b0;
    assign data[14300] = ~16'b0;
    assign data[14301] = ~16'b0;
    assign data[14302] = ~16'b0;
    assign data[14303] = ~16'b0;
    assign data[14304] = ~16'b0;
    assign data[14305] = ~16'b0;
    assign data[14306] = ~16'b0;
    assign data[14307] = ~16'b0;
    assign data[14308] = ~16'b0;
    assign data[14309] = ~16'b0;
    assign data[14310] = ~16'b0;
    assign data[14311] = ~16'b0;
    assign data[14312] = ~16'b0;
    assign data[14313] = ~16'b0;
    assign data[14314] = ~16'b0;
    assign data[14315] = ~16'b0;
    assign data[14316] = ~16'b0;
    assign data[14317] = ~16'b0;
    assign data[14318] = ~16'b0;
    assign data[14319] = ~16'b0;
    assign data[14320] = ~16'b0;
    assign data[14321] = ~16'b0;
    assign data[14322] = ~16'b0;
    assign data[14323] = ~16'b0;
    assign data[14324] = ~16'b0;
    assign data[14325] = ~16'b0;
    assign data[14326] = ~16'b0;
    assign data[14327] = ~16'b0;
    assign data[14328] = ~16'b0;
    assign data[14329] = ~16'b0;
    assign data[14330] = ~16'b0;
    assign data[14331] = ~16'b0;
    assign data[14332] = ~16'b0;
    assign data[14333] = ~16'b0;
    assign data[14334] = ~16'b0;
    assign data[14335] = ~16'b0;
    assign data[14336] = ~16'b0;
    assign data[14337] = ~16'b0;
    assign data[14338] = ~16'b0;
    assign data[14339] = ~16'b0;
    assign data[14340] = ~16'b0;
    assign data[14341] = ~16'b0;
    assign data[14342] = ~16'b0;
    assign data[14343] = ~16'b0;
    assign data[14344] = ~16'b0;
    assign data[14345] = ~16'b0;
    assign data[14346] = ~16'b0;
    assign data[14347] = ~16'b0;
    assign data[14348] = ~16'b0;
    assign data[14349] = ~16'b0;
    assign data[14350] = ~16'b0;
    assign data[14351] = ~16'b0;
    assign data[14352] = ~16'b0;
    assign data[14353] = ~16'b0;
    assign data[14354] = ~16'b0;
    assign data[14355] = ~16'b0;
    assign data[14356] = ~16'b0;
    assign data[14357] = ~16'b0;
    assign data[14358] = ~16'b0;
    assign data[14359] = ~16'b0;
    assign data[14360] = ~16'b0;
    assign data[14361] = ~16'b0;
    assign data[14362] = ~16'b0;
    assign data[14363] = ~16'b0;
    assign data[14364] = ~16'b0;
    assign data[14365] = ~16'b0;
    assign data[14366] = ~16'b0;
    assign data[14367] = ~16'b0;
    assign data[14368] = ~16'b0;
    assign data[14369] = ~16'b0;
    assign data[14370] = ~16'b0;
    assign data[14371] = ~16'b0;
    assign data[14372] = ~16'b0;
    assign data[14373] = ~16'b0;
    assign data[14374] = ~16'b0;
    assign data[14375] = ~16'b0;
    assign data[14376] = ~16'b0;
    assign data[14377] = ~16'b0;
    assign data[14378] = ~16'b0;
    assign data[14379] = ~16'b0;
    assign data[14380] = ~16'b0;
    assign data[14381] = ~16'b0;
    assign data[14382] = ~16'b0;
    assign data[14383] = ~16'b0;
    assign data[14384] = ~16'b0;
    assign data[14385] = ~16'b0;
    assign data[14386] = ~16'b0;
    assign data[14387] = ~16'b0;
    assign data[14388] = ~16'b0;
    assign data[14389] = ~16'b0;
    assign data[14390] = ~16'b0;
    assign data[14391] = ~16'b0;
    assign data[14392] = ~16'b0;
    assign data[14393] = ~16'b0;
    assign data[14394] = ~16'b0;
    assign data[14395] = ~16'b0;
    assign data[14396] = ~16'b0;
    assign data[14397] = ~16'b0;
    assign data[14398] = ~16'b0;
    assign data[14399] = ~16'b0;
    assign data[14400] = ~16'b0;
    assign data[14401] = ~16'b0;
    assign data[14402] = ~16'b0;
    assign data[14403] = ~16'b0;
    assign data[14404] = ~16'b0;
    assign data[14405] = ~16'b0;
    assign data[14406] = ~16'b0;
    assign data[14407] = ~16'b0;
    assign data[14408] = ~16'b0;
    assign data[14409] = ~16'b0;
    assign data[14410] = ~16'b0;
    assign data[14411] = ~16'b0;
    assign data[14412] = ~16'b0;
    assign data[14413] = ~16'b0;
    assign data[14414] = ~16'b0;
    assign data[14415] = ~16'b0;
    assign data[14416] = ~16'b0;
    assign data[14417] = ~16'b0;
    assign data[14418] = ~16'b0;
    assign data[14419] = ~16'b0;
    assign data[14420] = ~16'b0;
    assign data[14421] = ~16'b0;
    assign data[14422] = ~16'b0;
    assign data[14423] = ~16'b0;
    assign data[14424] = ~16'b0;
    assign data[14425] = ~16'b0;
    assign data[14426] = ~16'b0;
    assign data[14427] = ~16'b0;
    assign data[14428] = ~16'b0;
    assign data[14429] = ~16'b0;
    assign data[14430] = ~16'b0;
    assign data[14431] = ~16'b0;
    assign data[14432] = ~16'b0;
    assign data[14433] = ~16'b0;
    assign data[14434] = ~16'b0;
    assign data[14435] = ~16'b0;
    assign data[14436] = ~16'b0;
    assign data[14437] = ~16'b0;
    assign data[14438] = ~16'b0;
    assign data[14439] = ~16'b0;
    assign data[14440] = ~16'b0;
    assign data[14441] = ~16'b0;
    assign data[14442] = ~16'b0;
    assign data[14443] = ~16'b0;
    assign data[14444] = ~16'b0;
    assign data[14445] = ~16'b0;
    assign data[14446] = ~16'b0;
    assign data[14447] = ~16'b0;
    assign data[14448] = ~16'b0;
    assign data[14449] = ~16'b0;
    assign data[14450] = ~16'b0;
    assign data[14451] = ~16'b0;
    assign data[14452] = ~16'b0;
    assign data[14453] = ~16'b0;
    assign data[14454] = ~16'b0;
    assign data[14455] = ~16'b0;
    assign data[14456] = ~16'b0;
    assign data[14457] = ~16'b0;
    assign data[14458] = ~16'b0;
    assign data[14459] = ~16'b0;
    assign data[14460] = ~16'b0;
    assign data[14461] = ~16'b0;
    assign data[14462] = ~16'b0;
    assign data[14463] = ~16'b0;
    assign data[14464] = ~16'b0;
    assign data[14465] = ~16'b0;
    assign data[14466] = ~16'b0;
    assign data[14467] = ~16'b0;
    assign data[14468] = ~16'b0;
    assign data[14469] = ~16'b0;
    assign data[14470] = ~16'b0;
    assign data[14471] = ~16'b0;
    assign data[14472] = ~16'b0;
    assign data[14473] = ~16'b0;
    assign data[14474] = ~16'b0;
    assign data[14475] = ~16'b0;
    assign data[14476] = ~16'b0;
    assign data[14477] = ~16'b0;
    assign data[14478] = ~16'b0;
    assign data[14479] = ~16'b0;
    assign data[14480] = ~16'b0;
    assign data[14481] = ~16'b0;
    assign data[14482] = ~16'b0;
    assign data[14483] = ~16'b0;
    assign data[14484] = ~16'b0;
    assign data[14485] = ~16'b0;
    assign data[14486] = ~16'b0;
    assign data[14487] = ~16'b0;
    assign data[14488] = ~16'b0;
    assign data[14489] = ~16'b0;
    assign data[14490] = ~16'b0;
    assign data[14491] = ~16'b0;
    assign data[14492] = ~16'b0;
    assign data[14493] = ~16'b0;
    assign data[14494] = ~16'b0;
    assign data[14495] = ~16'b0;
    assign data[14496] = ~16'b0;
    assign data[14497] = ~16'b0;
    assign data[14498] = ~16'b0;
    assign data[14499] = ~16'b0;
    assign data[14500] = ~16'b0;
    assign data[14501] = ~16'b0;
    assign data[14502] = ~16'b0;
    assign data[14503] = ~16'b0;
    assign data[14504] = ~16'b0;
    assign data[14505] = ~16'b0;
    assign data[14506] = ~16'b0;
    assign data[14507] = ~16'b0;
    assign data[14508] = ~16'b0;
    assign data[14509] = ~16'b0;
    assign data[14510] = ~16'b0;
    assign data[14511] = ~16'b0;
    assign data[14512] = ~16'b0;
    assign data[14513] = ~16'b0;
    assign data[14514] = ~16'b0;
    assign data[14515] = ~16'b0;
    assign data[14516] = ~16'b0;
    assign data[14517] = ~16'b0;
    assign data[14518] = ~16'b0;
    assign data[14519] = ~16'b0;
    assign data[14520] = ~16'b0;
    assign data[14521] = ~16'b0;
    assign data[14522] = ~16'b0;
    assign data[14523] = ~16'b0;
    assign data[14524] = ~16'b0;
    assign data[14525] = ~16'b0;
    assign data[14526] = ~16'b0;
    assign data[14527] = ~16'b0;
    assign data[14528] = ~16'b0;
    assign data[14529] = ~16'b0;
    assign data[14530] = ~16'b0;
    assign data[14531] = ~16'b0;
    assign data[14532] = ~16'b0;
    assign data[14533] = ~16'b0;
    assign data[14534] = ~16'b0;
    assign data[14535] = ~16'b0;
    assign data[14536] = ~16'b0;
    assign data[14537] = ~16'b0;
    assign data[14538] = ~16'b0;
    assign data[14539] = ~16'b0;
    assign data[14540] = ~16'b0;
    assign data[14541] = ~16'b0;
    assign data[14542] = ~16'b0;
    assign data[14543] = ~16'b0;
    assign data[14544] = ~16'b0;
    assign data[14545] = ~16'b0;
    assign data[14546] = ~16'b0;
    assign data[14547] = ~16'b0;
    assign data[14548] = ~16'b0;
    assign data[14549] = ~16'b0;
    assign data[14550] = ~16'b0;
    assign data[14551] = ~16'b0;
    assign data[14552] = ~16'b0;
    assign data[14553] = ~16'b0;
    assign data[14554] = ~16'b0;
    assign data[14555] = ~16'b0;
    assign data[14556] = ~16'b0;
    assign data[14557] = ~16'b0;
    assign data[14558] = ~16'b0;
    assign data[14559] = ~16'b0;
    assign data[14560] = ~16'b0;
    assign data[14561] = ~16'b0;
    assign data[14562] = ~16'b0;
    assign data[14563] = ~16'b0;
    assign data[14564] = ~16'b0;
    assign data[14565] = ~16'b0;
    assign data[14566] = ~16'b0;
    assign data[14567] = ~16'b0;
    assign data[14568] = ~16'b0;
    assign data[14569] = ~16'b0;
    assign data[14570] = ~16'b0;
    assign data[14571] = ~16'b0;
    assign data[14572] = ~16'b0;
    assign data[14573] = ~16'b0;
    assign data[14574] = ~16'b0;
    assign data[14575] = ~16'b0;
    assign data[14576] = ~16'b0;
    assign data[14577] = ~16'b0;
    assign data[14578] = ~16'b0;
    assign data[14579] = ~16'b0;
    assign data[14580] = ~16'b0;
    assign data[14581] = ~16'b0;
    assign data[14582] = ~16'b0;
    assign data[14583] = ~16'b0;
    assign data[14584] = ~16'b0;
    assign data[14585] = ~16'b0;
    assign data[14586] = ~16'b0;
    assign data[14587] = ~16'b0;
    assign data[14588] = ~16'b0;
    assign data[14589] = ~16'b0;
    assign data[14590] = ~16'b0;
    assign data[14591] = ~16'b0;
    assign data[14592] = ~16'b0;
    assign data[14593] = ~16'b0;
    assign data[14594] = ~16'b0;
    assign data[14595] = ~16'b0;
    assign data[14596] = ~16'b0;
    assign data[14597] = ~16'b0;
    assign data[14598] = ~16'b0;
    assign data[14599] = ~16'b0;
    assign data[14600] = ~16'b0;
    assign data[14601] = ~16'b0;
    assign data[14602] = ~16'b0;
    assign data[14603] = ~16'b0;
    assign data[14604] = ~16'b0;
    assign data[14605] = ~16'b0;
    assign data[14606] = ~16'b0;
    assign data[14607] = ~16'b0;
    assign data[14608] = ~16'b0;
    assign data[14609] = ~16'b0;
    assign data[14610] = ~16'b0;
    assign data[14611] = ~16'b0;
    assign data[14612] = ~16'b0;
    assign data[14613] = ~16'b0;
    assign data[14614] = ~16'b0;
    assign data[14615] = ~16'b0;
    assign data[14616] = ~16'b0;
    assign data[14617] = ~16'b0;
    assign data[14618] = ~16'b0;
    assign data[14619] = ~16'b0;
    assign data[14620] = ~16'b0;
    assign data[14621] = ~16'b0;
    assign data[14622] = ~16'b0;
    assign data[14623] = ~16'b0;
    assign data[14624] = ~16'b0;
    assign data[14625] = ~16'b0;
    assign data[14626] = ~16'b0;
    assign data[14627] = ~16'b0;
    assign data[14628] = ~16'b0;
    assign data[14629] = ~16'b0;
    assign data[14630] = ~16'b0;
    assign data[14631] = ~16'b0;
    assign data[14632] = ~16'b0;
    assign data[14633] = ~16'b0;
    assign data[14634] = ~16'b0;
    assign data[14635] = ~16'b0;
    assign data[14636] = ~16'b0;
    assign data[14637] = ~16'b0;
    assign data[14638] = ~16'b0;
    assign data[14639] = ~16'b0;
    assign data[14640] = ~16'b0;
    assign data[14641] = ~16'b0;
    assign data[14642] = ~16'b0;
    assign data[14643] = ~16'b0;
    assign data[14644] = ~16'b0;
    assign data[14645] = ~16'b0;
    assign data[14646] = ~16'b0;
    assign data[14647] = ~16'b0;
    assign data[14648] = ~16'b0;
    assign data[14649] = ~16'b0;
    assign data[14650] = ~16'b0;
    assign data[14651] = ~16'b0;
    assign data[14652] = ~16'b0;
    assign data[14653] = ~16'b0;
    assign data[14654] = ~16'b0;
    assign data[14655] = ~16'b0;
    assign data[14656] = ~16'b0;
    assign data[14657] = ~16'b0;
    assign data[14658] = ~16'b0;
    assign data[14659] = ~16'b0;
    assign data[14660] = ~16'b0;
    assign data[14661] = ~16'b0;
    assign data[14662] = ~16'b0;
    assign data[14663] = ~16'b0;
    assign data[14664] = ~16'b0;
    assign data[14665] = ~16'b0;
    assign data[14666] = ~16'b0;
    assign data[14667] = ~16'b0;
    assign data[14668] = ~16'b0;
    assign data[14669] = ~16'b0;
    assign data[14670] = ~16'b0;
    assign data[14671] = ~16'b0;
    assign data[14672] = ~16'b0;
    assign data[14673] = ~16'b0;
    assign data[14674] = ~16'b0;
    assign data[14675] = ~16'b0;
    assign data[14676] = ~16'b0;
    assign data[14677] = ~16'b0;
    assign data[14678] = ~16'b0;
    assign data[14679] = ~16'b0;
    assign data[14680] = ~16'b0;
    assign data[14681] = ~16'b0;
    assign data[14682] = ~16'b0;
    assign data[14683] = ~16'b0;
    assign data[14684] = ~16'b0;
    assign data[14685] = ~16'b0;
    assign data[14686] = ~16'b0;
    assign data[14687] = ~16'b0;
    assign data[14688] = ~16'b0;
    assign data[14689] = ~16'b0;
    assign data[14690] = ~16'b0;
    assign data[14691] = ~16'b0;
    assign data[14692] = ~16'b0;
    assign data[14693] = ~16'b0;
    assign data[14694] = ~16'b0;
    assign data[14695] = ~16'b0;
    assign data[14696] = ~16'b0;
    assign data[14697] = ~16'b0;
    assign data[14698] = ~16'b0;
    assign data[14699] = ~16'b0;
    assign data[14700] = ~16'b0;
    assign data[14701] = ~16'b0;
    assign data[14702] = ~16'b0;
    assign data[14703] = ~16'b0;
    assign data[14704] = ~16'b0;
    assign data[14705] = ~16'b0;
    assign data[14706] = ~16'b0;
    assign data[14707] = ~16'b0;
    assign data[14708] = ~16'b0;
    assign data[14709] = ~16'b0;
    assign data[14710] = ~16'b0;
    assign data[14711] = ~16'b0;
    assign data[14712] = ~16'b0;
    assign data[14713] = ~16'b0;
    assign data[14714] = ~16'b0;
    assign data[14715] = ~16'b0;
    assign data[14716] = ~16'b0;
    assign data[14717] = ~16'b0;
    assign data[14718] = ~16'b0;
    assign data[14719] = ~16'b0;
    assign data[14720] = ~16'b0;
    assign data[14721] = ~16'b0;
    assign data[14722] = ~16'b0;
    assign data[14723] = ~16'b0;
    assign data[14724] = ~16'b0;
    assign data[14725] = ~16'b0;
    assign data[14726] = ~16'b0;
    assign data[14727] = ~16'b0;
    assign data[14728] = ~16'b0;
    assign data[14729] = ~16'b0;
    assign data[14730] = ~16'b0;
    assign data[14731] = ~16'b0;
    assign data[14732] = ~16'b0;
    assign data[14733] = ~16'b0;
    assign data[14734] = ~16'b0;
    assign data[14735] = ~16'b0;
    assign data[14736] = ~16'b0;
    assign data[14737] = ~16'b0;
    assign data[14738] = ~16'b0;
    assign data[14739] = ~16'b0;
    assign data[14740] = ~16'b0;
    assign data[14741] = ~16'b0;
    assign data[14742] = ~16'b0;
    assign data[14743] = ~16'b0;
    assign data[14744] = ~16'b0;
    assign data[14745] = ~16'b0;
    assign data[14746] = ~16'b0;
    assign data[14747] = ~16'b0;
    assign data[14748] = ~16'b0;
    assign data[14749] = ~16'b0;
    assign data[14750] = ~16'b0;
    assign data[14751] = ~16'b0;
    assign data[14752] = ~16'b0;
    assign data[14753] = ~16'b0;
    assign data[14754] = ~16'b0;
    assign data[14755] = ~16'b0;
    assign data[14756] = ~16'b0;
    assign data[14757] = ~16'b0;
    assign data[14758] = ~16'b0;
    assign data[14759] = ~16'b0;
    assign data[14760] = ~16'b0;
    assign data[14761] = ~16'b0;
    assign data[14762] = ~16'b0;
    assign data[14763] = ~16'b0;
    assign data[14764] = ~16'b0;
    assign data[14765] = ~16'b0;
    assign data[14766] = ~16'b0;
    assign data[14767] = ~16'b0;
    assign data[14768] = ~16'b0;
    assign data[14769] = ~16'b0;
    assign data[14770] = ~16'b0;
    assign data[14771] = ~16'b0;
    assign data[14772] = ~16'b0;
    assign data[14773] = ~16'b0;
    assign data[14774] = ~16'b0;
    assign data[14775] = ~16'b0;
    assign data[14776] = ~16'b0;
    assign data[14777] = ~16'b0;
    assign data[14778] = ~16'b0;
    assign data[14779] = ~16'b0;
    assign data[14780] = ~16'b0;
    assign data[14781] = ~16'b0;
    assign data[14782] = ~16'b0;
    assign data[14783] = ~16'b0;
    assign data[14784] = ~16'b0;
    assign data[14785] = ~16'b0;
    assign data[14786] = ~16'b0;
    assign data[14787] = ~16'b0;
    assign data[14788] = ~16'b0;
    assign data[14789] = ~16'b0;
    assign data[14790] = ~16'b0;
    assign data[14791] = ~16'b0;
    assign data[14792] = ~16'b0;
    assign data[14793] = ~16'b0;
    assign data[14794] = ~16'b0;
    assign data[14795] = ~16'b0;
    assign data[14796] = ~16'b0;
    assign data[14797] = ~16'b0;
    assign data[14798] = ~16'b0;
    assign data[14799] = ~16'b0;
    assign data[14800] = ~16'b0;
    assign data[14801] = ~16'b0;
    assign data[14802] = ~16'b0;
    assign data[14803] = ~16'b0;
    assign data[14804] = ~16'b0;
    assign data[14805] = ~16'b0;
    assign data[14806] = ~16'b0;
    assign data[14807] = ~16'b0;
    assign data[14808] = ~16'b0;
    assign data[14809] = ~16'b0;
    assign data[14810] = ~16'b0;
    assign data[14811] = ~16'b0;
    assign data[14812] = ~16'b0;
    assign data[14813] = ~16'b0;
    assign data[14814] = ~16'b0;
    assign data[14815] = ~16'b0;
    assign data[14816] = ~16'b0;
    assign data[14817] = ~16'b0;
    assign data[14818] = ~16'b0;
    assign data[14819] = ~16'b0;
    assign data[14820] = ~16'b0;
    assign data[14821] = ~16'b0;
    assign data[14822] = ~16'b0;
    assign data[14823] = ~16'b0;
    assign data[14824] = ~16'b0;
    assign data[14825] = ~16'b0;
    assign data[14826] = ~16'b0;
    assign data[14827] = ~16'b0;
    assign data[14828] = ~16'b0;
    assign data[14829] = ~16'b0;
    assign data[14830] = ~16'b0;
    assign data[14831] = ~16'b0;
    assign data[14832] = ~16'b0;
    assign data[14833] = ~16'b0;
    assign data[14834] = ~16'b0;
    assign data[14835] = ~16'b0;
    assign data[14836] = ~16'b0;
    assign data[14837] = ~16'b0;
    assign data[14838] = ~16'b0;
    assign data[14839] = ~16'b0;
    assign data[14840] = ~16'b0;
    assign data[14841] = ~16'b0;
    assign data[14842] = ~16'b0;
    assign data[14843] = ~16'b0;
    assign data[14844] = ~16'b0;
    assign data[14845] = ~16'b0;
    assign data[14846] = ~16'b0;
    assign data[14847] = ~16'b0;
    assign data[14848] = ~16'b0;
    assign data[14849] = ~16'b0;
    assign data[14850] = ~16'b0;
    assign data[14851] = ~16'b0;
    assign data[14852] = ~16'b0;
    assign data[14853] = ~16'b0;
    assign data[14854] = ~16'b0;
    assign data[14855] = ~16'b0;
    assign data[14856] = ~16'b0;
    assign data[14857] = ~16'b0;
    assign data[14858] = ~16'b0;
    assign data[14859] = ~16'b0;
    assign data[14860] = ~16'b0;
    assign data[14861] = ~16'b0;
    assign data[14862] = ~16'b0;
    assign data[14863] = ~16'b0;
    assign data[14864] = ~16'b0;
    assign data[14865] = ~16'b0;
    assign data[14866] = ~16'b0;
    assign data[14867] = ~16'b0;
    assign data[14868] = ~16'b0;
    assign data[14869] = ~16'b0;
    assign data[14870] = ~16'b0;
    assign data[14871] = ~16'b0;
    assign data[14872] = ~16'b0;
    assign data[14873] = ~16'b0;
    assign data[14874] = ~16'b0;
    assign data[14875] = ~16'b0;
    assign data[14876] = ~16'b0;
    assign data[14877] = ~16'b0;
    assign data[14878] = ~16'b0;
    assign data[14879] = ~16'b0;
    assign data[14880] = ~16'b0;
    assign data[14881] = ~16'b0;
    assign data[14882] = ~16'b0;
    assign data[14883] = ~16'b0;
    assign data[14884] = ~16'b0;
    assign data[14885] = ~16'b0;
    assign data[14886] = ~16'b0;
    assign data[14887] = ~16'b0;
    assign data[14888] = ~16'b0;
    assign data[14889] = ~16'b0;
    assign data[14890] = ~16'b0;
    assign data[14891] = ~16'b0;
    assign data[14892] = ~16'b0;
    assign data[14893] = ~16'b0;
    assign data[14894] = ~16'b0;
    assign data[14895] = ~16'b0;
    assign data[14896] = ~16'b0;
    assign data[14897] = ~16'b0;
    assign data[14898] = ~16'b0;
    assign data[14899] = ~16'b0;
    assign data[14900] = ~16'b0;
    assign data[14901] = ~16'b0;
    assign data[14902] = ~16'b0;
    assign data[14903] = ~16'b0;
    assign data[14904] = ~16'b0;
    assign data[14905] = ~16'b0;
    assign data[14906] = ~16'b0;
    assign data[14907] = ~16'b0;
    assign data[14908] = ~16'b0;
    assign data[14909] = ~16'b0;
    assign data[14910] = ~16'b0;
    assign data[14911] = ~16'b0;
    assign data[14912] = ~16'b0;
    assign data[14913] = ~16'b0;
    assign data[14914] = ~16'b0;
    assign data[14915] = ~16'b0;
    assign data[14916] = ~16'b0;
    assign data[14917] = ~16'b0;
    assign data[14918] = ~16'b0;
    assign data[14919] = ~16'b0;
    assign data[14920] = ~16'b0;
    assign data[14921] = ~16'b0;
    assign data[14922] = ~16'b0;
    assign data[14923] = ~16'b0;
    assign data[14924] = ~16'b0;
    assign data[14925] = ~16'b0;
    assign data[14926] = ~16'b0;
    assign data[14927] = ~16'b0;
    assign data[14928] = ~16'b0;
    assign data[14929] = ~16'b0;
    assign data[14930] = ~16'b0;
    assign data[14931] = ~16'b0;
    assign data[14932] = ~16'b0;
    assign data[14933] = ~16'b0;
    assign data[14934] = ~16'b0;
    assign data[14935] = ~16'b0;
    assign data[14936] = ~16'b0;
    assign data[14937] = ~16'b0;
    assign data[14938] = ~16'b0;
    assign data[14939] = ~16'b0;
    assign data[14940] = ~16'b0;
    assign data[14941] = ~16'b0;
    assign data[14942] = ~16'b0;
    assign data[14943] = ~16'b0;
    assign data[14944] = ~16'b0;
    assign data[14945] = ~16'b0;
    assign data[14946] = ~16'b0;
    assign data[14947] = ~16'b0;
    assign data[14948] = ~16'b0;
    assign data[14949] = ~16'b0;
    assign data[14950] = ~16'b0;
    assign data[14951] = ~16'b0;
    assign data[14952] = ~16'b0;
    assign data[14953] = ~16'b0;
    assign data[14954] = ~16'b0;
    assign data[14955] = ~16'b0;
    assign data[14956] = ~16'b0;
    assign data[14957] = ~16'b0;
    assign data[14958] = ~16'b0;
    assign data[14959] = ~16'b0;
    assign data[14960] = ~16'b0;
    assign data[14961] = ~16'b0;
    assign data[14962] = ~16'b0;
    assign data[14963] = ~16'b0;
    assign data[14964] = ~16'b0;
    assign data[14965] = ~16'b0;
    assign data[14966] = ~16'b0;
    assign data[14967] = ~16'b0;
    assign data[14968] = ~16'b0;
    assign data[14969] = ~16'b0;
    assign data[14970] = ~16'b0;
    assign data[14971] = ~16'b0;
    assign data[14972] = ~16'b0;
    assign data[14973] = ~16'b0;
    assign data[14974] = ~16'b0;
    assign data[14975] = ~16'b0;
    assign data[14976] = ~16'b0;
    assign data[14977] = ~16'b0;
    assign data[14978] = ~16'b0;
    assign data[14979] = ~16'b0;
    assign data[14980] = ~16'b0;
    assign data[14981] = ~16'b0;
    assign data[14982] = ~16'b0;
    assign data[14983] = ~16'b0;
    assign data[14984] = ~16'b0;
    assign data[14985] = ~16'b0;
    assign data[14986] = ~16'b0;
    assign data[14987] = ~16'b0;
    assign data[14988] = ~16'b0;
    assign data[14989] = ~16'b0;
    assign data[14990] = ~16'b0;
    assign data[14991] = ~16'b0;
    assign data[14992] = ~16'b0;
    assign data[14993] = ~16'b0;
    assign data[14994] = ~16'b0;
    assign data[14995] = ~16'b0;
    assign data[14996] = ~16'b0;
    assign data[14997] = ~16'b0;
    assign data[14998] = ~16'b0;
    assign data[14999] = ~16'b0;
    assign data[15000] = ~16'b0;
    assign data[15001] = ~16'b0;
    assign data[15002] = ~16'b0;
    assign data[15003] = ~16'b0;
    assign data[15004] = ~16'b0;
    assign data[15005] = ~16'b0;
    assign data[15006] = ~16'b0;
    assign data[15007] = ~16'b0;
    assign data[15008] = ~16'b0;
    assign data[15009] = ~16'b0;
    assign data[15010] = ~16'b0;
    assign data[15011] = ~16'b0;
    assign data[15012] = ~16'b0;
    assign data[15013] = ~16'b0;
    assign data[15014] = ~16'b0;
    assign data[15015] = ~16'b0;
    assign data[15016] = ~16'b0;
    assign data[15017] = ~16'b0;
    assign data[15018] = ~16'b0;
    assign data[15019] = ~16'b0;
endmodule


