`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/25/2023 05:03:22 PM
// Design Name: 
// Module Name: audio_game_oled
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module audio_game_oled(
    input clock, clk_os, clk_display, clk_pos,
    input [10:0] num, 
    input [6:0] x,y,
    output [15:0] oled_data
    );
    
    parameter reg gravity = 5;
    reg flag = 0;
    reg [4:0] y_acc;
    wire [4:0] y_acceleration;
    wire x_move;
    wire [31:0] offset;
    wire [1:0] stop_x;
    always @ (posedge clock) begin
        if (num >= 0 && num < 205)
            begin  
                y_acc <= 0;
                flag <= 0;
            end
        else if (num >= 205 && num < 409)
            begin
                y_acc <= 50;
                flag <= 1;
            end
        else if (num >= 409 && num < 614)
            begin
                y_acc <= 45;
                flag <= 1;            
            end
        else if (num >= 614 && num < 819)
            begin
                y_acc <= 40;
                flag <= 1;            
            end
        else if (num >= 819 && num < 1024)
            begin 
                y_acc <= 35;
                flag <= 1;            
            end
        else if (num >= 1024 && num < 1229)
            begin 
                y_acc <= 30;
                flag <= 1;            
            end
        else if (num >= 1229 && num < 1434)
            begin
                y_acc <= 25;
                flag <= 1;            
            end
        else if (num >= 1434 && num < 1638)
            begin
                y_acc <= 20;
                flag <= 1;            
            end
        else if (num >= 1638 && num < 1842)
            begin
                y_acc <= 15;
                flag <= 1;            
            end
        else if (num >= 1842 && num <= 2047)
            begin 
                y_acc <= 10;
                flag <= 1;            
            end
    end
    
    assign y_acceleration = y_acc;
    assign x_move = flag && stop_x;
    
    check_x_offset x_offset(clk_os, x_move, offset);
    output_display oled(clk_display, clk_pos, y_acceleration, x,y,offset, stop_x, oled_data);
endmodule


module check_x_offset(
    input clk10Hz, x_move,
    output reg [31:0] offset = 0
);

    parameter max_offset = 642;
    always @ (posedge clk10Hz) begin
        if (x_move) begin
            offset <= (offset == max_offset) ? 0 : offset + 1;
        end
    end
    
endmodule

module output_display(
    input clk_display, clk_pos,
    input [4:0] y_acc,
    input [6:0] x,y,
    input [31:0] offset,
    output reg [1:0] stop_x = 1,
    output reg [15:0] oled_data
);

    wire [15:0] data [0:7379];
    wire [31:0] index;
    assign index = (x * 10) + (y - 54) + (10 * offset);
    
    parameter square_size = 3;
    parameter max_y_speed = 10;
    parameter max_y_pos = 3;
    parameter min_y_pos = 60;
    
    wire square_pos;
    //initial position of ball
    reg [6:0] x_pos = 31;
    reg [6:0] y_pos = 20; 
    
    reg [31:0] count = 0;
    
    // boolean logics 
    wire hit_top, hit_bottom, hit_right, on_land;
    wire index_to_check_right;
    wire [31:0] index_to_check_bottom [0:6];
    
    //death screen
    wire [15:0] death_oled;
    
    //assign all boolean logic here
    assign hit_top = (y_pos <= max_y_pos);
    assign hit_bottom = (y_pos >= min_y_pos);
    assign index_to_check_right = 350 + (y_pos + square_size - 54) + 10 * offset;
    assign index_to_check_bottom[0] = 280 + offset * 10;
    assign index_to_check_bottom[1] = 290 + offset * 10;
    assign index_to_check_bottom[2] = 300 + offset * 10;
    assign index_to_check_bottom[3] = 310 + offset * 10;
    assign index_to_check_bottom[4] = 320 + offset * 10;
    assign index_to_check_bottom[5] = 330 + offset * 10;
    assign index_to_check_bottom[6] = 340 + offset * 10;
    assign hit_right = (y_pos > 50) && (data[index_to_check_right] == 16'b0);
    assign on_land = (y_pos == 50) && (data[index_to_check_bottom[0]] == 16'b0 || 
                                       data[index_to_check_bottom[1]] == 16'b0 || 
                                       data[index_to_check_bottom[2]] == 16'b0 || 
                                       data[index_to_check_bottom[3]] == 16'b0 || 
                                       data[index_to_check_bottom[4]] == 16'b0 || 
                                       data[index_to_check_bottom[5]] == 16'b0 || 
                                       data[index_to_check_bottom[6]] == 16'b0);
    
    //output logic of x,y coordinates to render the square
    assign square_pos  = (x >= x_pos - square_size && x <= x_pos + square_size) &&
                         (y >= y_pos - square_size && y <= y_pos + square_size);
                         
                        
    always @(posedge clk_display) begin
        stop_x <= hit_right || hit_bottom ? 0 : 1;
        oled_data <= hit_bottom ? death_oled : square_pos ? 16'b0 : y > 53 ? data[index] : ~16'b0;
    end
    
    always @(posedge clk_pos) begin
        //y_speed = (y_speed >= max_y_speed) && (y_acc > 0) ? max_y_speed : y_speed + y_acc;
        if (y_acc > 0) begin
            count <= count >= y_acc - 1 ? 0 : count + 1;
            y_pos <= count == y_acc - 1? (hit_top ? max_y_pos : hit_bottom ? min_y_pos : y_pos - 1) : y_pos;
        end
        
        else begin
            count <= count >= 34 ? 0 : count + 1;
            y_pos <= count == 34 ? (hit_bottom ? min_y_pos : on_land ? 50 : y_pos + 1) : y_pos;
        end
    end
    
    
    death_image d1(.x(x), .y(y), .oled_data(death_oled));
    
    assign data[0] = 16'b0;
    assign data[1] = 16'b0;
    assign data[2] = 16'b0;
    assign data[3] = 16'b0;
    assign data[4] = 16'b0;
    assign data[5] = 16'b0;
    assign data[6] = 16'b0;
    assign data[7] = 16'b0;
    assign data[8] = 16'b0;
    assign data[9] = 16'b0;
    assign data[10] = 16'b0;
    assign data[11] = 16'b0;
    assign data[12] = 16'b0;
    assign data[13] = 16'b0;
    assign data[14] = 16'b0;
    assign data[15] = 16'b0;
    assign data[16] = 16'b0;
    assign data[17] = 16'b0;
    assign data[18] = 16'b0;
    assign data[19] = 16'b0;
    assign data[20] = 16'b0;
    assign data[21] = 16'b0;
    assign data[22] = ~16'b0;
    assign data[23] = ~16'b0;
    assign data[24] = ~16'b0;
    assign data[25] = ~16'b0;
    assign data[26] = ~16'b0;
    assign data[27] = ~16'b0;
    assign data[28] = ~16'b0;
    assign data[29] = ~16'b0;
    assign data[30] = 16'b0;
    assign data[31] = 16'b0;
    assign data[32] = ~16'b0;
    assign data[33] = ~16'b0;
    assign data[34] = ~16'b0;
    assign data[35] = ~16'b0;
    assign data[36] = ~16'b0;
    assign data[37] = ~16'b0;
    assign data[38] = ~16'b0;
    assign data[39] = ~16'b0;
    assign data[40] = 16'b0;
    assign data[41] = 16'b0;
    assign data[42] = ~16'b0;
    assign data[43] = ~16'b0;
    assign data[44] = ~16'b0;
    assign data[45] = ~16'b0;
    assign data[46] = ~16'b0;
    assign data[47] = ~16'b0;
    assign data[48] = ~16'b0;
    assign data[49] = ~16'b0;
    assign data[50] = 16'b0;
    assign data[51] = 16'b0;
    assign data[52] = ~16'b0;
    assign data[53] = ~16'b0;
    assign data[54] = ~16'b0;
    assign data[55] = ~16'b0;
    assign data[56] = ~16'b0;
    assign data[57] = ~16'b0;
    assign data[58] = ~16'b0;
    assign data[59] = ~16'b0;
    assign data[60] = 16'b0;
    assign data[61] = 16'b0;
    assign data[62] = ~16'b0;
    assign data[63] = ~16'b0;
    assign data[64] = ~16'b0;
    assign data[65] = ~16'b0;
    assign data[66] = ~16'b0;
    assign data[67] = ~16'b0;
    assign data[68] = ~16'b0;
    assign data[69] = ~16'b0;
    assign data[70] = 16'b0;
    assign data[71] = 16'b0;
    assign data[72] = ~16'b0;
    assign data[73] = ~16'b0;
    assign data[74] = ~16'b0;
    assign data[75] = ~16'b0;
    assign data[76] = ~16'b0;
    assign data[77] = ~16'b0;
    assign data[78] = ~16'b0;
    assign data[79] = ~16'b0;
    assign data[80] = 16'b0;
    assign data[81] = 16'b0;
    assign data[82] = ~16'b0;
    assign data[83] = ~16'b0;
    assign data[84] = ~16'b0;
    assign data[85] = ~16'b0;
    assign data[86] = ~16'b0;
    assign data[87] = ~16'b0;
    assign data[88] = ~16'b0;
    assign data[89] = ~16'b0;
    assign data[90] = 16'b0;
    assign data[91] = 16'b0;
    assign data[92] = ~16'b0;
    assign data[93] = ~16'b0;
    assign data[94] = ~16'b0;
    assign data[95] = ~16'b0;
    assign data[96] = ~16'b0;
    assign data[97] = ~16'b0;
    assign data[98] = ~16'b0;
    assign data[99] = ~16'b0;
    assign data[100] = 16'b0;
    assign data[101] = 16'b0;
    assign data[102] = ~16'b0;
    assign data[103] = ~16'b0;
    assign data[104] = ~16'b0;
    assign data[105] = ~16'b0;
    assign data[106] = ~16'b0;
    assign data[107] = ~16'b0;
    assign data[108] = ~16'b0;
    assign data[109] = ~16'b0;
    assign data[110] = 16'b0;
    assign data[111] = 16'b0;
    assign data[112] = ~16'b0;
    assign data[113] = ~16'b0;
    assign data[114] = ~16'b0;
    assign data[115] = ~16'b0;
    assign data[116] = ~16'b0;
    assign data[117] = ~16'b0;
    assign data[118] = ~16'b0;
    assign data[119] = ~16'b0;
    assign data[120] = 16'b0;
    assign data[121] = 16'b0;
    assign data[122] = ~16'b0;
    assign data[123] = ~16'b0;
    assign data[124] = ~16'b0;
    assign data[125] = ~16'b0;
    assign data[126] = ~16'b0;
    assign data[127] = ~16'b0;
    assign data[128] = ~16'b0;
    assign data[129] = ~16'b0;
    assign data[130] = 16'b0;
    assign data[131] = 16'b0;
    assign data[132] = ~16'b0;
    assign data[133] = ~16'b0;
    assign data[134] = ~16'b0;
    assign data[135] = ~16'b0;
    assign data[136] = ~16'b0;
    assign data[137] = ~16'b0;
    assign data[138] = ~16'b0;
    assign data[139] = ~16'b0;
    assign data[140] = 16'b0;
    assign data[141] = 16'b0;
    assign data[142] = ~16'b0;
    assign data[143] = ~16'b0;
    assign data[144] = ~16'b0;
    assign data[145] = ~16'b0;
    assign data[146] = ~16'b0;
    assign data[147] = ~16'b0;
    assign data[148] = ~16'b0;
    assign data[149] = ~16'b0;
    assign data[150] = 16'b0;
    assign data[151] = 16'b0;
    assign data[152] = ~16'b0;
    assign data[153] = ~16'b0;
    assign data[154] = ~16'b0;
    assign data[155] = ~16'b0;
    assign data[156] = ~16'b0;
    assign data[157] = ~16'b0;
    assign data[158] = ~16'b0;
    assign data[159] = ~16'b0;
    assign data[160] = 16'b0;
    assign data[161] = 16'b0;
    assign data[162] = ~16'b0;
    assign data[163] = ~16'b0;
    assign data[164] = ~16'b0;
    assign data[165] = ~16'b0;
    assign data[166] = ~16'b0;
    assign data[167] = ~16'b0;
    assign data[168] = ~16'b0;
    assign data[169] = ~16'b0;
    assign data[170] = 16'b0;
    assign data[171] = 16'b0;
    assign data[172] = ~16'b0;
    assign data[173] = ~16'b0;
    assign data[174] = ~16'b0;
    assign data[175] = ~16'b0;
    assign data[176] = ~16'b0;
    assign data[177] = ~16'b0;
    assign data[178] = ~16'b0;
    assign data[179] = ~16'b0;
    assign data[180] = 16'b0;
    assign data[181] = 16'b0;
    assign data[182] = ~16'b0;
    assign data[183] = ~16'b0;
    assign data[184] = ~16'b0;
    assign data[185] = ~16'b0;
    assign data[186] = ~16'b0;
    assign data[187] = ~16'b0;
    assign data[188] = ~16'b0;
    assign data[189] = ~16'b0;
    assign data[190] = 16'b0;
    assign data[191] = 16'b0;
    assign data[192] = ~16'b0;
    assign data[193] = ~16'b0;
    assign data[194] = ~16'b0;
    assign data[195] = ~16'b0;
    assign data[196] = ~16'b0;
    assign data[197] = ~16'b0;
    assign data[198] = ~16'b0;
    assign data[199] = ~16'b0;
    assign data[200] = 16'b0;
    assign data[201] = 16'b0;
    assign data[202] = ~16'b0;
    assign data[203] = ~16'b0;
    assign data[204] = ~16'b0;
    assign data[205] = ~16'b0;
    assign data[206] = ~16'b0;
    assign data[207] = ~16'b0;
    assign data[208] = ~16'b0;
    assign data[209] = ~16'b0;
    assign data[210] = 16'b0;
    assign data[211] = 16'b0;
    assign data[212] = ~16'b0;
    assign data[213] = ~16'b0;
    assign data[214] = ~16'b0;
    assign data[215] = ~16'b0;
    assign data[216] = ~16'b0;
    assign data[217] = ~16'b0;
    assign data[218] = ~16'b0;
    assign data[219] = ~16'b0;
    assign data[220] = 16'b0;
    assign data[221] = 16'b0;
    assign data[222] = ~16'b0;
    assign data[223] = ~16'b0;
    assign data[224] = ~16'b0;
    assign data[225] = ~16'b0;
    assign data[226] = ~16'b0;
    assign data[227] = ~16'b0;
    assign data[228] = ~16'b0;
    assign data[229] = ~16'b0;
    assign data[230] = 16'b0;
    assign data[231] = 16'b0;
    assign data[232] = ~16'b0;
    assign data[233] = ~16'b0;
    assign data[234] = ~16'b0;
    assign data[235] = ~16'b0;
    assign data[236] = ~16'b0;
    assign data[237] = ~16'b0;
    assign data[238] = ~16'b0;
    assign data[239] = ~16'b0;
    assign data[240] = 16'b0;
    assign data[241] = 16'b0;
    assign data[242] = ~16'b0;
    assign data[243] = ~16'b0;
    assign data[244] = ~16'b0;
    assign data[245] = ~16'b0;
    assign data[246] = ~16'b0;
    assign data[247] = ~16'b0;
    assign data[248] = ~16'b0;
    assign data[249] = ~16'b0;
    assign data[250] = 16'b0;
    assign data[251] = 16'b0;
    assign data[252] = ~16'b0;
    assign data[253] = ~16'b0;
    assign data[254] = ~16'b0;
    assign data[255] = ~16'b0;
    assign data[256] = ~16'b0;
    assign data[257] = ~16'b0;
    assign data[258] = ~16'b0;
    assign data[259] = ~16'b0;
    assign data[260] = 16'b0;
    assign data[261] = 16'b0;
    assign data[262] = ~16'b0;
    assign data[263] = ~16'b0;
    assign data[264] = ~16'b0;
    assign data[265] = ~16'b0;
    assign data[266] = ~16'b0;
    assign data[267] = ~16'b0;
    assign data[268] = ~16'b0;
    assign data[269] = ~16'b0;
    assign data[270] = 16'b0;
    assign data[271] = 16'b0;
    assign data[272] = ~16'b0;
    assign data[273] = ~16'b0;
    assign data[274] = ~16'b0;
    assign data[275] = ~16'b0;
    assign data[276] = ~16'b0;
    assign data[277] = ~16'b0;
    assign data[278] = ~16'b0;
    assign data[279] = ~16'b0;
    assign data[280] = 16'b0;
    assign data[281] = 16'b0;
    assign data[282] = ~16'b0;
    assign data[283] = ~16'b0;
    assign data[284] = ~16'b0;
    assign data[285] = ~16'b0;
    assign data[286] = ~16'b0;
    assign data[287] = ~16'b0;
    assign data[288] = ~16'b0;
    assign data[289] = ~16'b0;
    assign data[290] = 16'b0;
    assign data[291] = 16'b0;
    assign data[292] = ~16'b0;
    assign data[293] = ~16'b0;
    assign data[294] = ~16'b0;
    assign data[295] = ~16'b0;
    assign data[296] = ~16'b0;
    assign data[297] = ~16'b0;
    assign data[298] = ~16'b0;
    assign data[299] = ~16'b0;
    assign data[300] = 16'b0;
    assign data[301] = 16'b0;
    assign data[302] = ~16'b0;
    assign data[303] = ~16'b0;
    assign data[304] = ~16'b0;
    assign data[305] = ~16'b0;
    assign data[306] = ~16'b0;
    assign data[307] = ~16'b0;
    assign data[308] = ~16'b0;
    assign data[309] = ~16'b0;
    assign data[310] = 16'b0;
    assign data[311] = 16'b0;
    assign data[312] = ~16'b0;
    assign data[313] = ~16'b0;
    assign data[314] = ~16'b0;
    assign data[315] = ~16'b0;
    assign data[316] = ~16'b0;
    assign data[317] = ~16'b0;
    assign data[318] = ~16'b0;
    assign data[319] = ~16'b0;
    assign data[320] = 16'b0;
    assign data[321] = 16'b0;
    assign data[322] = ~16'b0;
    assign data[323] = ~16'b0;
    assign data[324] = ~16'b0;
    assign data[325] = ~16'b0;
    assign data[326] = ~16'b0;
    assign data[327] = ~16'b0;
    assign data[328] = ~16'b0;
    assign data[329] = ~16'b0;
    assign data[330] = 16'b0;
    assign data[331] = 16'b0;
    assign data[332] = ~16'b0;
    assign data[333] = ~16'b0;
    assign data[334] = ~16'b0;
    assign data[335] = ~16'b0;
    assign data[336] = ~16'b0;
    assign data[337] = ~16'b0;
    assign data[338] = ~16'b0;
    assign data[339] = ~16'b0;
    assign data[340] = 16'b0;
    assign data[341] = 16'b0;
    assign data[342] = ~16'b0;
    assign data[343] = ~16'b0;
    assign data[344] = ~16'b0;
    assign data[345] = ~16'b0;
    assign data[346] = ~16'b0;
    assign data[347] = ~16'b0;
    assign data[348] = ~16'b0;
    assign data[349] = ~16'b0;
    assign data[350] = 16'b0;
    assign data[351] = 16'b0;
    assign data[352] = ~16'b0;
    assign data[353] = ~16'b0;
    assign data[354] = ~16'b0;
    assign data[355] = ~16'b0;
    assign data[356] = ~16'b0;
    assign data[357] = ~16'b0;
    assign data[358] = ~16'b0;
    assign data[359] = ~16'b0;
    assign data[360] = 16'b0;
    assign data[361] = 16'b0;
    assign data[362] = ~16'b0;
    assign data[363] = ~16'b0;
    assign data[364] = ~16'b0;
    assign data[365] = ~16'b0;
    assign data[366] = ~16'b0;
    assign data[367] = ~16'b0;
    assign data[368] = ~16'b0;
    assign data[369] = ~16'b0;
    assign data[370] = 16'b0;
    assign data[371] = 16'b0;
    assign data[372] = ~16'b0;
    assign data[373] = ~16'b0;
    assign data[374] = ~16'b0;
    assign data[375] = ~16'b0;
    assign data[376] = ~16'b0;
    assign data[377] = ~16'b0;
    assign data[378] = ~16'b0;
    assign data[379] = ~16'b0;
    assign data[380] = 16'b0;
    assign data[381] = 16'b0;
    assign data[382] = ~16'b0;
    assign data[383] = ~16'b0;
    assign data[384] = ~16'b0;
    assign data[385] = ~16'b0;
    assign data[386] = ~16'b0;
    assign data[387] = ~16'b0;
    assign data[388] = ~16'b0;
    assign data[389] = ~16'b0;
    assign data[390] = 16'b0;
    assign data[391] = 16'b0;
    assign data[392] = ~16'b0;
    assign data[393] = ~16'b0;
    assign data[394] = ~16'b0;
    assign data[395] = ~16'b0;
    assign data[396] = ~16'b0;
    assign data[397] = ~16'b0;
    assign data[398] = ~16'b0;
    assign data[399] = ~16'b0;
    assign data[400] = 16'b0;
    assign data[401] = 16'b0;
    assign data[402] = ~16'b0;
    assign data[403] = ~16'b0;
    assign data[404] = ~16'b0;
    assign data[405] = ~16'b0;
    assign data[406] = ~16'b0;
    assign data[407] = ~16'b0;
    assign data[408] = ~16'b0;
    assign data[409] = ~16'b0;
    assign data[410] = 16'b0;
    assign data[411] = 16'b0;
    assign data[412] = ~16'b0;
    assign data[413] = ~16'b0;
    assign data[414] = ~16'b0;
    assign data[415] = ~16'b0;
    assign data[416] = ~16'b0;
    assign data[417] = ~16'b0;
    assign data[418] = ~16'b0;
    assign data[419] = ~16'b0;
    assign data[420] = 16'b0;
    assign data[421] = 16'b0;
    assign data[422] = ~16'b0;
    assign data[423] = ~16'b0;
    assign data[424] = ~16'b0;
    assign data[425] = ~16'b0;
    assign data[426] = ~16'b0;
    assign data[427] = ~16'b0;
    assign data[428] = ~16'b0;
    assign data[429] = ~16'b0;
    assign data[430] = 16'b0;
    assign data[431] = 16'b0;
    assign data[432] = ~16'b0;
    assign data[433] = ~16'b0;
    assign data[434] = ~16'b0;
    assign data[435] = ~16'b0;
    assign data[436] = ~16'b0;
    assign data[437] = ~16'b0;
    assign data[438] = ~16'b0;
    assign data[439] = ~16'b0;
    assign data[440] = 16'b0;
    assign data[441] = 16'b0;
    assign data[442] = ~16'b0;
    assign data[443] = ~16'b0;
    assign data[444] = ~16'b0;
    assign data[445] = ~16'b0;
    assign data[446] = ~16'b0;
    assign data[447] = ~16'b0;
    assign data[448] = ~16'b0;
    assign data[449] = ~16'b0;
    assign data[450] = 16'b0;
    assign data[451] = 16'b0;
    assign data[452] = ~16'b0;
    assign data[453] = ~16'b0;
    assign data[454] = ~16'b0;
    assign data[455] = ~16'b0;
    assign data[456] = ~16'b0;
    assign data[457] = ~16'b0;
    assign data[458] = ~16'b0;
    assign data[459] = ~16'b0;
    assign data[460] = 16'b0;
    assign data[461] = 16'b0;
    assign data[462] = ~16'b0;
    assign data[463] = ~16'b0;
    assign data[464] = ~16'b0;
    assign data[465] = ~16'b0;
    assign data[466] = ~16'b0;
    assign data[467] = ~16'b0;
    assign data[468] = ~16'b0;
    assign data[469] = ~16'b0;
    assign data[470] = 16'b0;
    assign data[471] = 16'b0;
    assign data[472] = ~16'b0;
    assign data[473] = ~16'b0;
    assign data[474] = ~16'b0;
    assign data[475] = ~16'b0;
    assign data[476] = ~16'b0;
    assign data[477] = ~16'b0;
    assign data[478] = ~16'b0;
    assign data[479] = ~16'b0;
    assign data[480] = 16'b0;
    assign data[481] = 16'b0;
    assign data[482] = ~16'b0;
    assign data[483] = ~16'b0;
    assign data[484] = ~16'b0;
    assign data[485] = ~16'b0;
    assign data[486] = ~16'b0;
    assign data[487] = ~16'b0;
    assign data[488] = ~16'b0;
    assign data[489] = ~16'b0;
    assign data[490] = 16'b0;
    assign data[491] = 16'b0;
    assign data[492] = ~16'b0;
    assign data[493] = ~16'b0;
    assign data[494] = ~16'b0;
    assign data[495] = ~16'b0;
    assign data[496] = ~16'b0;
    assign data[497] = ~16'b0;
    assign data[498] = ~16'b0;
    assign data[499] = ~16'b0;
    assign data[500] = 16'b0;
    assign data[501] = 16'b0;
    assign data[502] = ~16'b0;
    assign data[503] = ~16'b0;
    assign data[504] = ~16'b0;
    assign data[505] = ~16'b0;
    assign data[506] = ~16'b0;
    assign data[507] = ~16'b0;
    assign data[508] = ~16'b0;
    assign data[509] = ~16'b0;
    assign data[510] = 16'b0;
    assign data[511] = 16'b0;
    assign data[512] = ~16'b0;
    assign data[513] = ~16'b0;
    assign data[514] = ~16'b0;
    assign data[515] = ~16'b0;
    assign data[516] = ~16'b0;
    assign data[517] = ~16'b0;
    assign data[518] = ~16'b0;
    assign data[519] = ~16'b0;
    assign data[520] = 16'b0;
    assign data[521] = 16'b0;
    assign data[522] = ~16'b0;
    assign data[523] = ~16'b0;
    assign data[524] = ~16'b0;
    assign data[525] = ~16'b0;
    assign data[526] = ~16'b0;
    assign data[527] = ~16'b0;
    assign data[528] = ~16'b0;
    assign data[529] = ~16'b0;
    assign data[530] = 16'b0;
    assign data[531] = 16'b0;
    assign data[532] = ~16'b0;
    assign data[533] = ~16'b0;
    assign data[534] = ~16'b0;
    assign data[535] = ~16'b0;
    assign data[536] = ~16'b0;
    assign data[537] = ~16'b0;
    assign data[538] = ~16'b0;
    assign data[539] = ~16'b0;
    assign data[540] = 16'b0;
    assign data[541] = 16'b0;
    assign data[542] = 16'b0;
    assign data[543] = 16'b0;
    assign data[544] = 16'b0;
    assign data[545] = 16'b0;
    assign data[546] = 16'b0;
    assign data[547] = 16'b0;
    assign data[548] = 16'b0;
    assign data[549] = 16'b0;
    assign data[550] = 16'b0;
    assign data[551] = 16'b0;
    assign data[552] = 16'b0;
    assign data[553] = 16'b0;
    assign data[554] = 16'b0;
    assign data[555] = 16'b0;
    assign data[556] = 16'b0;
    assign data[557] = 16'b0;
    assign data[558] = 16'b0;
    assign data[559] = 16'b0;
    assign data[560] = ~16'b0;
    assign data[561] = ~16'b0;
    assign data[562] = ~16'b0;
    assign data[563] = ~16'b0;
    assign data[564] = ~16'b0;
    assign data[565] = ~16'b0;
    assign data[566] = ~16'b0;
    assign data[567] = ~16'b0;
    assign data[568] = ~16'b0;
    assign data[569] = ~16'b0;
    assign data[570] = ~16'b0;
    assign data[571] = ~16'b0;
    assign data[572] = ~16'b0;
    assign data[573] = ~16'b0;
    assign data[574] = ~16'b0;
    assign data[575] = ~16'b0;
    assign data[576] = ~16'b0;
    assign data[577] = ~16'b0;
    assign data[578] = ~16'b0;
    assign data[579] = ~16'b0;
    assign data[580] = ~16'b0;
    assign data[581] = ~16'b0;
    assign data[582] = ~16'b0;
    assign data[583] = ~16'b0;
    assign data[584] = ~16'b0;
    assign data[585] = ~16'b0;
    assign data[586] = ~16'b0;
    assign data[587] = ~16'b0;
    assign data[588] = ~16'b0;
    assign data[589] = ~16'b0;
    assign data[590] = ~16'b0;
    assign data[591] = ~16'b0;
    assign data[592] = ~16'b0;
    assign data[593] = ~16'b0;
    assign data[594] = ~16'b0;
    assign data[595] = ~16'b0;
    assign data[596] = ~16'b0;
    assign data[597] = ~16'b0;
    assign data[598] = ~16'b0;
    assign data[599] = ~16'b0;
    assign data[600] = ~16'b0;
    assign data[601] = ~16'b0;
    assign data[602] = ~16'b0;
    assign data[603] = ~16'b0;
    assign data[604] = ~16'b0;
    assign data[605] = ~16'b0;
    assign data[606] = ~16'b0;
    assign data[607] = ~16'b0;
    assign data[608] = ~16'b0;
    assign data[609] = ~16'b0;
    assign data[610] = ~16'b0;
    assign data[611] = ~16'b0;
    assign data[612] = ~16'b0;
    assign data[613] = ~16'b0;
    assign data[614] = ~16'b0;
    assign data[615] = ~16'b0;
    assign data[616] = ~16'b0;
    assign data[617] = ~16'b0;
    assign data[618] = ~16'b0;
    assign data[619] = ~16'b0;
    assign data[620] = ~16'b0;
    assign data[621] = ~16'b0;
    assign data[622] = ~16'b0;
    assign data[623] = ~16'b0;
    assign data[624] = ~16'b0;
    assign data[625] = ~16'b0;
    assign data[626] = ~16'b0;
    assign data[627] = ~16'b0;
    assign data[628] = ~16'b0;
    assign data[629] = ~16'b0;
    assign data[630] = ~16'b0;
    assign data[631] = ~16'b0;
    assign data[632] = ~16'b0;
    assign data[633] = ~16'b0;
    assign data[634] = ~16'b0;
    assign data[635] = ~16'b0;
    assign data[636] = ~16'b0;
    assign data[637] = ~16'b0;
    assign data[638] = ~16'b0;
    assign data[639] = ~16'b0;
    assign data[640] = ~16'b0;
    assign data[641] = ~16'b0;
    assign data[642] = ~16'b0;
    assign data[643] = ~16'b0;
    assign data[644] = ~16'b0;
    assign data[645] = ~16'b0;
    assign data[646] = ~16'b0;
    assign data[647] = ~16'b0;
    assign data[648] = ~16'b0;
    assign data[649] = ~16'b0;
    assign data[650] = ~16'b0;
    assign data[651] = ~16'b0;
    assign data[652] = ~16'b0;
    assign data[653] = ~16'b0;
    assign data[654] = ~16'b0;
    assign data[655] = ~16'b0;
    assign data[656] = ~16'b0;
    assign data[657] = ~16'b0;
    assign data[658] = ~16'b0;
    assign data[659] = ~16'b0;
    assign data[660] = ~16'b0;
    assign data[661] = ~16'b0;
    assign data[662] = ~16'b0;
    assign data[663] = ~16'b0;
    assign data[664] = ~16'b0;
    assign data[665] = ~16'b0;
    assign data[666] = ~16'b0;
    assign data[667] = ~16'b0;
    assign data[668] = ~16'b0;
    assign data[669] = ~16'b0;
    assign data[670] = ~16'b0;
    assign data[671] = ~16'b0;
    assign data[672] = ~16'b0;
    assign data[673] = ~16'b0;
    assign data[674] = ~16'b0;
    assign data[675] = ~16'b0;
    assign data[676] = ~16'b0;
    assign data[677] = ~16'b0;
    assign data[678] = ~16'b0;
    assign data[679] = ~16'b0;
    assign data[680] = ~16'b0;
    assign data[681] = ~16'b0;
    assign data[682] = ~16'b0;
    assign data[683] = ~16'b0;
    assign data[684] = ~16'b0;
    assign data[685] = ~16'b0;
    assign data[686] = ~16'b0;
    assign data[687] = ~16'b0;
    assign data[688] = ~16'b0;
    assign data[689] = ~16'b0;
    assign data[690] = ~16'b0;
    assign data[691] = ~16'b0;
    assign data[692] = ~16'b0;
    assign data[693] = ~16'b0;
    assign data[694] = ~16'b0;
    assign data[695] = ~16'b0;
    assign data[696] = ~16'b0;
    assign data[697] = ~16'b0;
    assign data[698] = ~16'b0;
    assign data[699] = ~16'b0;
    assign data[700] = ~16'b0;
    assign data[701] = ~16'b0;
    assign data[702] = ~16'b0;
    assign data[703] = ~16'b0;
    assign data[704] = ~16'b0;
    assign data[705] = ~16'b0;
    assign data[706] = ~16'b0;
    assign data[707] = ~16'b0;
    assign data[708] = ~16'b0;
    assign data[709] = ~16'b0;
    assign data[710] = ~16'b0;
    assign data[711] = ~16'b0;
    assign data[712] = ~16'b0;
    assign data[713] = ~16'b0;
    assign data[714] = ~16'b0;
    assign data[715] = ~16'b0;
    assign data[716] = ~16'b0;
    assign data[717] = ~16'b0;
    assign data[718] = ~16'b0;
    assign data[719] = ~16'b0;
    assign data[720] = ~16'b0;
    assign data[721] = ~16'b0;
    assign data[722] = ~16'b0;
    assign data[723] = ~16'b0;
    assign data[724] = ~16'b0;
    assign data[725] = ~16'b0;
    assign data[726] = ~16'b0;
    assign data[727] = ~16'b0;
    assign data[728] = ~16'b0;
    assign data[729] = ~16'b0;
    assign data[730] = ~16'b0;
    assign data[731] = ~16'b0;
    assign data[732] = ~16'b0;
    assign data[733] = ~16'b0;
    assign data[734] = ~16'b0;
    assign data[735] = ~16'b0;
    assign data[736] = ~16'b0;
    assign data[737] = ~16'b0;
    assign data[738] = ~16'b0;
    assign data[739] = ~16'b0;
    assign data[740] = ~16'b0;
    assign data[741] = ~16'b0;
    assign data[742] = ~16'b0;
    assign data[743] = ~16'b0;
    assign data[744] = ~16'b0;
    assign data[745] = ~16'b0;
    assign data[746] = ~16'b0;
    assign data[747] = ~16'b0;
    assign data[748] = ~16'b0;
    assign data[749] = ~16'b0;
    assign data[750] = ~16'b0;
    assign data[751] = ~16'b0;
    assign data[752] = ~16'b0;
    assign data[753] = ~16'b0;
    assign data[754] = ~16'b0;
    assign data[755] = ~16'b0;
    assign data[756] = ~16'b0;
    assign data[757] = ~16'b0;
    assign data[758] = ~16'b0;
    assign data[759] = ~16'b0;
    assign data[760] = 16'b0;
    assign data[761] = 16'b0;
    assign data[762] = 16'b0;
    assign data[763] = 16'b0;
    assign data[764] = 16'b0;
    assign data[765] = 16'b0;
    assign data[766] = 16'b0;
    assign data[767] = 16'b0;
    assign data[768] = 16'b0;
    assign data[769] = 16'b0;
    assign data[770] = 16'b0;
    assign data[771] = 16'b0;
    assign data[772] = 16'b0;
    assign data[773] = 16'b0;
    assign data[774] = 16'b0;
    assign data[775] = 16'b0;
    assign data[776] = 16'b0;
    assign data[777] = 16'b0;
    assign data[778] = 16'b0;
    assign data[779] = 16'b0;
    assign data[780] = 16'b0;
    assign data[781] = 16'b0;
    assign data[782] = ~16'b0;
    assign data[783] = ~16'b0;
    assign data[784] = ~16'b0;
    assign data[785] = ~16'b0;
    assign data[786] = ~16'b0;
    assign data[787] = ~16'b0;
    assign data[788] = ~16'b0;
    assign data[789] = ~16'b0;
    assign data[790] = 16'b0;
    assign data[791] = 16'b0;
    assign data[792] = ~16'b0;
    assign data[793] = ~16'b0;
    assign data[794] = ~16'b0;
    assign data[795] = ~16'b0;
    assign data[796] = ~16'b0;
    assign data[797] = ~16'b0;
    assign data[798] = ~16'b0;
    assign data[799] = ~16'b0;
    assign data[800] = 16'b0;
    assign data[801] = 16'b0;
    assign data[802] = ~16'b0;
    assign data[803] = ~16'b0;
    assign data[804] = ~16'b0;
    assign data[805] = ~16'b0;
    assign data[806] = ~16'b0;
    assign data[807] = ~16'b0;
    assign data[808] = ~16'b0;
    assign data[809] = ~16'b0;
    assign data[810] = 16'b0;
    assign data[811] = 16'b0;
    assign data[812] = ~16'b0;
    assign data[813] = ~16'b0;
    assign data[814] = ~16'b0;
    assign data[815] = ~16'b0;
    assign data[816] = ~16'b0;
    assign data[817] = ~16'b0;
    assign data[818] = ~16'b0;
    assign data[819] = ~16'b0;
    assign data[820] = 16'b0;
    assign data[821] = 16'b0;
    assign data[822] = ~16'b0;
    assign data[823] = ~16'b0;
    assign data[824] = ~16'b0;
    assign data[825] = ~16'b0;
    assign data[826] = ~16'b0;
    assign data[827] = ~16'b0;
    assign data[828] = ~16'b0;
    assign data[829] = ~16'b0;
    assign data[830] = 16'b0;
    assign data[831] = 16'b0;
    assign data[832] = ~16'b0;
    assign data[833] = ~16'b0;
    assign data[834] = ~16'b0;
    assign data[835] = ~16'b0;
    assign data[836] = ~16'b0;
    assign data[837] = ~16'b0;
    assign data[838] = ~16'b0;
    assign data[839] = ~16'b0;
    assign data[840] = 16'b0;
    assign data[841] = 16'b0;
    assign data[842] = ~16'b0;
    assign data[843] = ~16'b0;
    assign data[844] = ~16'b0;
    assign data[845] = ~16'b0;
    assign data[846] = ~16'b0;
    assign data[847] = ~16'b0;
    assign data[848] = ~16'b0;
    assign data[849] = ~16'b0;
    assign data[850] = 16'b0;
    assign data[851] = 16'b0;
    assign data[852] = ~16'b0;
    assign data[853] = ~16'b0;
    assign data[854] = ~16'b0;
    assign data[855] = ~16'b0;
    assign data[856] = ~16'b0;
    assign data[857] = ~16'b0;
    assign data[858] = ~16'b0;
    assign data[859] = ~16'b0;
    assign data[860] = 16'b0;
    assign data[861] = 16'b0;
    assign data[862] = ~16'b0;
    assign data[863] = ~16'b0;
    assign data[864] = ~16'b0;
    assign data[865] = ~16'b0;
    assign data[866] = ~16'b0;
    assign data[867] = ~16'b0;
    assign data[868] = ~16'b0;
    assign data[869] = ~16'b0;
    assign data[870] = 16'b0;
    assign data[871] = 16'b0;
    assign data[872] = ~16'b0;
    assign data[873] = ~16'b0;
    assign data[874] = ~16'b0;
    assign data[875] = ~16'b0;
    assign data[876] = ~16'b0;
    assign data[877] = ~16'b0;
    assign data[878] = ~16'b0;
    assign data[879] = ~16'b0;
    assign data[880] = 16'b0;
    assign data[881] = 16'b0;
    assign data[882] = ~16'b0;
    assign data[883] = ~16'b0;
    assign data[884] = ~16'b0;
    assign data[885] = ~16'b0;
    assign data[886] = ~16'b0;
    assign data[887] = ~16'b0;
    assign data[888] = ~16'b0;
    assign data[889] = ~16'b0;
    assign data[890] = 16'b0;
    assign data[891] = 16'b0;
    assign data[892] = ~16'b0;
    assign data[893] = ~16'b0;
    assign data[894] = ~16'b0;
    assign data[895] = ~16'b0;
    assign data[896] = ~16'b0;
    assign data[897] = ~16'b0;
    assign data[898] = ~16'b0;
    assign data[899] = ~16'b0;
    assign data[900] = 16'b0;
    assign data[901] = 16'b0;
    assign data[902] = ~16'b0;
    assign data[903] = ~16'b0;
    assign data[904] = ~16'b0;
    assign data[905] = ~16'b0;
    assign data[906] = ~16'b0;
    assign data[907] = ~16'b0;
    assign data[908] = ~16'b0;
    assign data[909] = ~16'b0;
    assign data[910] = 16'b0;
    assign data[911] = 16'b0;
    assign data[912] = ~16'b0;
    assign data[913] = ~16'b0;
    assign data[914] = ~16'b0;
    assign data[915] = ~16'b0;
    assign data[916] = ~16'b0;
    assign data[917] = ~16'b0;
    assign data[918] = ~16'b0;
    assign data[919] = ~16'b0;
    assign data[920] = 16'b0;
    assign data[921] = 16'b0;
    assign data[922] = ~16'b0;
    assign data[923] = ~16'b0;
    assign data[924] = ~16'b0;
    assign data[925] = ~16'b0;
    assign data[926] = ~16'b0;
    assign data[927] = ~16'b0;
    assign data[928] = ~16'b0;
    assign data[929] = ~16'b0;
    assign data[930] = 16'b0;
    assign data[931] = 16'b0;
    assign data[932] = ~16'b0;
    assign data[933] = ~16'b0;
    assign data[934] = ~16'b0;
    assign data[935] = ~16'b0;
    assign data[936] = ~16'b0;
    assign data[937] = ~16'b0;
    assign data[938] = ~16'b0;
    assign data[939] = ~16'b0;
    assign data[940] = 16'b0;
    assign data[941] = 16'b0;
    assign data[942] = ~16'b0;
    assign data[943] = ~16'b0;
    assign data[944] = ~16'b0;
    assign data[945] = ~16'b0;
    assign data[946] = ~16'b0;
    assign data[947] = ~16'b0;
    assign data[948] = ~16'b0;
    assign data[949] = ~16'b0;
    assign data[950] = 16'b0;
    assign data[951] = 16'b0;
    assign data[952] = ~16'b0;
    assign data[953] = ~16'b0;
    assign data[954] = ~16'b0;
    assign data[955] = ~16'b0;
    assign data[956] = ~16'b0;
    assign data[957] = ~16'b0;
    assign data[958] = ~16'b0;
    assign data[959] = ~16'b0;
    assign data[960] = 16'b0;
    assign data[961] = 16'b0;
    assign data[962] = ~16'b0;
    assign data[963] = ~16'b0;
    assign data[964] = ~16'b0;
    assign data[965] = ~16'b0;
    assign data[966] = ~16'b0;
    assign data[967] = ~16'b0;
    assign data[968] = ~16'b0;
    assign data[969] = ~16'b0;
    assign data[970] = 16'b0;
    assign data[971] = 16'b0;
    assign data[972] = 16'b0;
    assign data[973] = 16'b0;
    assign data[974] = 16'b0;
    assign data[975] = 16'b0;
    assign data[976] = 16'b0;
    assign data[977] = 16'b0;
    assign data[978] = 16'b0;
    assign data[979] = 16'b0;
    assign data[980] = 16'b0;
    assign data[981] = 16'b0;
    assign data[982] = 16'b0;
    assign data[983] = 16'b0;
    assign data[984] = 16'b0;
    assign data[985] = 16'b0;
    assign data[986] = 16'b0;
    assign data[987] = 16'b0;
    assign data[988] = 16'b0;
    assign data[989] = 16'b0;
    assign data[990] = ~16'b0;
    assign data[991] = ~16'b0;
    assign data[992] = ~16'b0;
    assign data[993] = ~16'b0;
    assign data[994] = ~16'b0;
    assign data[995] = ~16'b0;
    assign data[996] = ~16'b0;
    assign data[997] = ~16'b0;
    assign data[998] = ~16'b0;
    assign data[999] = ~16'b0;
    assign data[1000] = ~16'b0;
    assign data[1001] = ~16'b0;
    assign data[1002] = ~16'b0;
    assign data[1003] = ~16'b0;
    assign data[1004] = ~16'b0;
    assign data[1005] = ~16'b0;
    assign data[1006] = ~16'b0;
    assign data[1007] = ~16'b0;
    assign data[1008] = ~16'b0;
    assign data[1009] = ~16'b0;
    assign data[1010] = ~16'b0;
    assign data[1011] = ~16'b0;
    assign data[1012] = ~16'b0;
    assign data[1013] = ~16'b0;
    assign data[1014] = ~16'b0;
    assign data[1015] = ~16'b0;
    assign data[1016] = ~16'b0;
    assign data[1017] = ~16'b0;
    assign data[1018] = ~16'b0;
    assign data[1019] = ~16'b0;
    assign data[1020] = ~16'b0;
    assign data[1021] = ~16'b0;
    assign data[1022] = ~16'b0;
    assign data[1023] = ~16'b0;
    assign data[1024] = ~16'b0;
    assign data[1025] = ~16'b0;
    assign data[1026] = ~16'b0;
    assign data[1027] = ~16'b0;
    assign data[1028] = ~16'b0;
    assign data[1029] = ~16'b0;
    assign data[1030] = ~16'b0;
    assign data[1031] = ~16'b0;
    assign data[1032] = ~16'b0;
    assign data[1033] = ~16'b0;
    assign data[1034] = ~16'b0;
    assign data[1035] = ~16'b0;
    assign data[1036] = ~16'b0;
    assign data[1037] = ~16'b0;
    assign data[1038] = ~16'b0;
    assign data[1039] = ~16'b0;
    assign data[1040] = ~16'b0;
    assign data[1041] = ~16'b0;
    assign data[1042] = ~16'b0;
    assign data[1043] = ~16'b0;
    assign data[1044] = ~16'b0;
    assign data[1045] = ~16'b0;
    assign data[1046] = ~16'b0;
    assign data[1047] = ~16'b0;
    assign data[1048] = ~16'b0;
    assign data[1049] = ~16'b0;
    assign data[1050] = ~16'b0;
    assign data[1051] = ~16'b0;
    assign data[1052] = ~16'b0;
    assign data[1053] = ~16'b0;
    assign data[1054] = ~16'b0;
    assign data[1055] = ~16'b0;
    assign data[1056] = ~16'b0;
    assign data[1057] = ~16'b0;
    assign data[1058] = ~16'b0;
    assign data[1059] = ~16'b0;
    assign data[1060] = ~16'b0;
    assign data[1061] = ~16'b0;
    assign data[1062] = ~16'b0;
    assign data[1063] = ~16'b0;
    assign data[1064] = ~16'b0;
    assign data[1065] = ~16'b0;
    assign data[1066] = ~16'b0;
    assign data[1067] = ~16'b0;
    assign data[1068] = ~16'b0;
    assign data[1069] = ~16'b0;
    assign data[1070] = ~16'b0;
    assign data[1071] = ~16'b0;
    assign data[1072] = ~16'b0;
    assign data[1073] = ~16'b0;
    assign data[1074] = ~16'b0;
    assign data[1075] = ~16'b0;
    assign data[1076] = ~16'b0;
    assign data[1077] = ~16'b0;
    assign data[1078] = ~16'b0;
    assign data[1079] = ~16'b0;
    assign data[1080] = ~16'b0;
    assign data[1081] = ~16'b0;
    assign data[1082] = ~16'b0;
    assign data[1083] = ~16'b0;
    assign data[1084] = ~16'b0;
    assign data[1085] = ~16'b0;
    assign data[1086] = ~16'b0;
    assign data[1087] = ~16'b0;
    assign data[1088] = ~16'b0;
    assign data[1089] = ~16'b0;
    assign data[1090] = ~16'b0;
    assign data[1091] = ~16'b0;
    assign data[1092] = ~16'b0;
    assign data[1093] = ~16'b0;
    assign data[1094] = ~16'b0;
    assign data[1095] = ~16'b0;
    assign data[1096] = ~16'b0;
    assign data[1097] = ~16'b0;
    assign data[1098] = ~16'b0;
    assign data[1099] = ~16'b0;
    assign data[1100] = ~16'b0;
    assign data[1101] = ~16'b0;
    assign data[1102] = ~16'b0;
    assign data[1103] = ~16'b0;
    assign data[1104] = ~16'b0;
    assign data[1105] = ~16'b0;
    assign data[1106] = ~16'b0;
    assign data[1107] = ~16'b0;
    assign data[1108] = ~16'b0;
    assign data[1109] = ~16'b0;
    assign data[1110] = ~16'b0;
    assign data[1111] = ~16'b0;
    assign data[1112] = ~16'b0;
    assign data[1113] = ~16'b0;
    assign data[1114] = ~16'b0;
    assign data[1115] = ~16'b0;
    assign data[1116] = ~16'b0;
    assign data[1117] = ~16'b0;
    assign data[1118] = ~16'b0;
    assign data[1119] = ~16'b0;
    assign data[1120] = ~16'b0;
    assign data[1121] = ~16'b0;
    assign data[1122] = ~16'b0;
    assign data[1123] = ~16'b0;
    assign data[1124] = ~16'b0;
    assign data[1125] = ~16'b0;
    assign data[1126] = ~16'b0;
    assign data[1127] = ~16'b0;
    assign data[1128] = ~16'b0;
    assign data[1129] = ~16'b0;
    assign data[1130] = ~16'b0;
    assign data[1131] = ~16'b0;
    assign data[1132] = ~16'b0;
    assign data[1133] = ~16'b0;
    assign data[1134] = ~16'b0;
    assign data[1135] = ~16'b0;
    assign data[1136] = ~16'b0;
    assign data[1137] = ~16'b0;
    assign data[1138] = ~16'b0;
    assign data[1139] = ~16'b0;
    assign data[1140] = ~16'b0;
    assign data[1141] = ~16'b0;
    assign data[1142] = ~16'b0;
    assign data[1143] = ~16'b0;
    assign data[1144] = ~16'b0;
    assign data[1145] = ~16'b0;
    assign data[1146] = ~16'b0;
    assign data[1147] = ~16'b0;
    assign data[1148] = ~16'b0;
    assign data[1149] = ~16'b0;
    assign data[1150] = ~16'b0;
    assign data[1151] = ~16'b0;
    assign data[1152] = ~16'b0;
    assign data[1153] = ~16'b0;
    assign data[1154] = ~16'b0;
    assign data[1155] = ~16'b0;
    assign data[1156] = ~16'b0;
    assign data[1157] = ~16'b0;
    assign data[1158] = ~16'b0;
    assign data[1159] = ~16'b0;
    assign data[1160] = ~16'b0;
    assign data[1161] = ~16'b0;
    assign data[1162] = ~16'b0;
    assign data[1163] = ~16'b0;
    assign data[1164] = ~16'b0;
    assign data[1165] = ~16'b0;
    assign data[1166] = ~16'b0;
    assign data[1167] = ~16'b0;
    assign data[1168] = ~16'b0;
    assign data[1169] = ~16'b0;
    assign data[1170] = ~16'b0;
    assign data[1171] = ~16'b0;
    assign data[1172] = ~16'b0;
    assign data[1173] = ~16'b0;
    assign data[1174] = ~16'b0;
    assign data[1175] = ~16'b0;
    assign data[1176] = ~16'b0;
    assign data[1177] = ~16'b0;
    assign data[1178] = ~16'b0;
    assign data[1179] = ~16'b0;
    assign data[1180] = ~16'b0;
    assign data[1181] = ~16'b0;
    assign data[1182] = ~16'b0;
    assign data[1183] = ~16'b0;
    assign data[1184] = ~16'b0;
    assign data[1185] = ~16'b0;
    assign data[1186] = ~16'b0;
    assign data[1187] = ~16'b0;
    assign data[1188] = ~16'b0;
    assign data[1189] = ~16'b0;
    assign data[1190] = ~16'b0;
    assign data[1191] = ~16'b0;
    assign data[1192] = ~16'b0;
    assign data[1193] = ~16'b0;
    assign data[1194] = ~16'b0;
    assign data[1195] = ~16'b0;
    assign data[1196] = ~16'b0;
    assign data[1197] = ~16'b0;
    assign data[1198] = ~16'b0;
    assign data[1199] = ~16'b0;
    assign data[1200] = 16'b0;
    assign data[1201] = 16'b0;
    assign data[1202] = 16'b0;
    assign data[1203] = 16'b0;
    assign data[1204] = 16'b0;
    assign data[1205] = 16'b0;
    assign data[1206] = 16'b0;
    assign data[1207] = 16'b0;
    assign data[1208] = 16'b0;
    assign data[1209] = 16'b0;
    assign data[1210] = 16'b0;
    assign data[1211] = 16'b0;
    assign data[1212] = 16'b0;
    assign data[1213] = 16'b0;
    assign data[1214] = 16'b0;
    assign data[1215] = 16'b0;
    assign data[1216] = 16'b0;
    assign data[1217] = 16'b0;
    assign data[1218] = 16'b0;
    assign data[1219] = 16'b0;
    assign data[1220] = 16'b0;
    assign data[1221] = 16'b0;
    assign data[1222] = ~16'b0;
    assign data[1223] = ~16'b0;
    assign data[1224] = ~16'b0;
    assign data[1225] = ~16'b0;
    assign data[1226] = ~16'b0;
    assign data[1227] = ~16'b0;
    assign data[1228] = ~16'b0;
    assign data[1229] = ~16'b0;
    assign data[1230] = 16'b0;
    assign data[1231] = 16'b0;
    assign data[1232] = ~16'b0;
    assign data[1233] = ~16'b0;
    assign data[1234] = ~16'b0;
    assign data[1235] = ~16'b0;
    assign data[1236] = ~16'b0;
    assign data[1237] = ~16'b0;
    assign data[1238] = ~16'b0;
    assign data[1239] = ~16'b0;
    assign data[1240] = 16'b0;
    assign data[1241] = 16'b0;
    assign data[1242] = ~16'b0;
    assign data[1243] = ~16'b0;
    assign data[1244] = ~16'b0;
    assign data[1245] = ~16'b0;
    assign data[1246] = ~16'b0;
    assign data[1247] = ~16'b0;
    assign data[1248] = ~16'b0;
    assign data[1249] = ~16'b0;
    assign data[1250] = 16'b0;
    assign data[1251] = 16'b0;
    assign data[1252] = ~16'b0;
    assign data[1253] = ~16'b0;
    assign data[1254] = ~16'b0;
    assign data[1255] = ~16'b0;
    assign data[1256] = ~16'b0;
    assign data[1257] = ~16'b0;
    assign data[1258] = ~16'b0;
    assign data[1259] = ~16'b0;
    assign data[1260] = 16'b0;
    assign data[1261] = 16'b0;
    assign data[1262] = ~16'b0;
    assign data[1263] = ~16'b0;
    assign data[1264] = ~16'b0;
    assign data[1265] = ~16'b0;
    assign data[1266] = ~16'b0;
    assign data[1267] = ~16'b0;
    assign data[1268] = ~16'b0;
    assign data[1269] = ~16'b0;
    assign data[1270] = 16'b0;
    assign data[1271] = 16'b0;
    assign data[1272] = ~16'b0;
    assign data[1273] = ~16'b0;
    assign data[1274] = ~16'b0;
    assign data[1275] = ~16'b0;
    assign data[1276] = ~16'b0;
    assign data[1277] = ~16'b0;
    assign data[1278] = ~16'b0;
    assign data[1279] = ~16'b0;
    assign data[1280] = 16'b0;
    assign data[1281] = 16'b0;
    assign data[1282] = ~16'b0;
    assign data[1283] = ~16'b0;
    assign data[1284] = ~16'b0;
    assign data[1285] = ~16'b0;
    assign data[1286] = ~16'b0;
    assign data[1287] = ~16'b0;
    assign data[1288] = ~16'b0;
    assign data[1289] = ~16'b0;
    assign data[1290] = 16'b0;
    assign data[1291] = 16'b0;
    assign data[1292] = ~16'b0;
    assign data[1293] = ~16'b0;
    assign data[1294] = ~16'b0;
    assign data[1295] = ~16'b0;
    assign data[1296] = ~16'b0;
    assign data[1297] = ~16'b0;
    assign data[1298] = ~16'b0;
    assign data[1299] = ~16'b0;
    assign data[1300] = 16'b0;
    assign data[1301] = 16'b0;
    assign data[1302] = ~16'b0;
    assign data[1303] = ~16'b0;
    assign data[1304] = ~16'b0;
    assign data[1305] = ~16'b0;
    assign data[1306] = ~16'b0;
    assign data[1307] = ~16'b0;
    assign data[1308] = ~16'b0;
    assign data[1309] = ~16'b0;
    assign data[1310] = 16'b0;
    assign data[1311] = 16'b0;
    assign data[1312] = ~16'b0;
    assign data[1313] = ~16'b0;
    assign data[1314] = ~16'b0;
    assign data[1315] = ~16'b0;
    assign data[1316] = ~16'b0;
    assign data[1317] = ~16'b0;
    assign data[1318] = ~16'b0;
    assign data[1319] = ~16'b0;
    assign data[1320] = 16'b0;
    assign data[1321] = 16'b0;
    assign data[1322] = ~16'b0;
    assign data[1323] = ~16'b0;
    assign data[1324] = ~16'b0;
    assign data[1325] = ~16'b0;
    assign data[1326] = ~16'b0;
    assign data[1327] = ~16'b0;
    assign data[1328] = ~16'b0;
    assign data[1329] = ~16'b0;
    assign data[1330] = 16'b0;
    assign data[1331] = 16'b0;
    assign data[1332] = ~16'b0;
    assign data[1333] = ~16'b0;
    assign data[1334] = ~16'b0;
    assign data[1335] = ~16'b0;
    assign data[1336] = ~16'b0;
    assign data[1337] = ~16'b0;
    assign data[1338] = ~16'b0;
    assign data[1339] = ~16'b0;
    assign data[1340] = 16'b0;
    assign data[1341] = 16'b0;
    assign data[1342] = ~16'b0;
    assign data[1343] = ~16'b0;
    assign data[1344] = ~16'b0;
    assign data[1345] = ~16'b0;
    assign data[1346] = ~16'b0;
    assign data[1347] = ~16'b0;
    assign data[1348] = ~16'b0;
    assign data[1349] = ~16'b0;
    assign data[1350] = 16'b0;
    assign data[1351] = 16'b0;
    assign data[1352] = ~16'b0;
    assign data[1353] = ~16'b0;
    assign data[1354] = ~16'b0;
    assign data[1355] = ~16'b0;
    assign data[1356] = ~16'b0;
    assign data[1357] = ~16'b0;
    assign data[1358] = ~16'b0;
    assign data[1359] = ~16'b0;
    assign data[1360] = 16'b0;
    assign data[1361] = 16'b0;
    assign data[1362] = ~16'b0;
    assign data[1363] = ~16'b0;
    assign data[1364] = ~16'b0;
    assign data[1365] = ~16'b0;
    assign data[1366] = ~16'b0;
    assign data[1367] = ~16'b0;
    assign data[1368] = ~16'b0;
    assign data[1369] = ~16'b0;
    assign data[1370] = 16'b0;
    assign data[1371] = 16'b0;
    assign data[1372] = ~16'b0;
    assign data[1373] = ~16'b0;
    assign data[1374] = ~16'b0;
    assign data[1375] = ~16'b0;
    assign data[1376] = ~16'b0;
    assign data[1377] = ~16'b0;
    assign data[1378] = ~16'b0;
    assign data[1379] = ~16'b0;
    assign data[1380] = 16'b0;
    assign data[1381] = 16'b0;
    assign data[1382] = ~16'b0;
    assign data[1383] = ~16'b0;
    assign data[1384] = ~16'b0;
    assign data[1385] = ~16'b0;
    assign data[1386] = ~16'b0;
    assign data[1387] = ~16'b0;
    assign data[1388] = ~16'b0;
    assign data[1389] = ~16'b0;
    assign data[1390] = 16'b0;
    assign data[1391] = 16'b0;
    assign data[1392] = ~16'b0;
    assign data[1393] = ~16'b0;
    assign data[1394] = ~16'b0;
    assign data[1395] = ~16'b0;
    assign data[1396] = ~16'b0;
    assign data[1397] = ~16'b0;
    assign data[1398] = ~16'b0;
    assign data[1399] = ~16'b0;
    assign data[1400] = 16'b0;
    assign data[1401] = 16'b0;
    assign data[1402] = ~16'b0;
    assign data[1403] = ~16'b0;
    assign data[1404] = ~16'b0;
    assign data[1405] = ~16'b0;
    assign data[1406] = ~16'b0;
    assign data[1407] = ~16'b0;
    assign data[1408] = ~16'b0;
    assign data[1409] = ~16'b0;
    assign data[1410] = 16'b0;
    assign data[1411] = 16'b0;
    assign data[1412] = ~16'b0;
    assign data[1413] = ~16'b0;
    assign data[1414] = ~16'b0;
    assign data[1415] = ~16'b0;
    assign data[1416] = ~16'b0;
    assign data[1417] = ~16'b0;
    assign data[1418] = ~16'b0;
    assign data[1419] = ~16'b0;
    assign data[1420] = 16'b0;
    assign data[1421] = 16'b0;
    assign data[1422] = ~16'b0;
    assign data[1423] = ~16'b0;
    assign data[1424] = ~16'b0;
    assign data[1425] = ~16'b0;
    assign data[1426] = ~16'b0;
    assign data[1427] = ~16'b0;
    assign data[1428] = ~16'b0;
    assign data[1429] = ~16'b0;
    assign data[1430] = 16'b0;
    assign data[1431] = 16'b0;
    assign data[1432] = ~16'b0;
    assign data[1433] = ~16'b0;
    assign data[1434] = ~16'b0;
    assign data[1435] = ~16'b0;
    assign data[1436] = ~16'b0;
    assign data[1437] = ~16'b0;
    assign data[1438] = ~16'b0;
    assign data[1439] = ~16'b0;
    assign data[1440] = 16'b0;
    assign data[1441] = 16'b0;
    assign data[1442] = ~16'b0;
    assign data[1443] = ~16'b0;
    assign data[1444] = ~16'b0;
    assign data[1445] = ~16'b0;
    assign data[1446] = ~16'b0;
    assign data[1447] = ~16'b0;
    assign data[1448] = ~16'b0;
    assign data[1449] = ~16'b0;
    assign data[1450] = 16'b0;
    assign data[1451] = 16'b0;
    assign data[1452] = ~16'b0;
    assign data[1453] = ~16'b0;
    assign data[1454] = ~16'b0;
    assign data[1455] = ~16'b0;
    assign data[1456] = ~16'b0;
    assign data[1457] = ~16'b0;
    assign data[1458] = ~16'b0;
    assign data[1459] = ~16'b0;
    assign data[1460] = 16'b0;
    assign data[1461] = 16'b0;
    assign data[1462] = ~16'b0;
    assign data[1463] = ~16'b0;
    assign data[1464] = ~16'b0;
    assign data[1465] = ~16'b0;
    assign data[1466] = ~16'b0;
    assign data[1467] = ~16'b0;
    assign data[1468] = ~16'b0;
    assign data[1469] = ~16'b0;
    assign data[1470] = 16'b0;
    assign data[1471] = 16'b0;
    assign data[1472] = ~16'b0;
    assign data[1473] = ~16'b0;
    assign data[1474] = ~16'b0;
    assign data[1475] = ~16'b0;
    assign data[1476] = ~16'b0;
    assign data[1477] = ~16'b0;
    assign data[1478] = ~16'b0;
    assign data[1479] = ~16'b0;
    assign data[1480] = 16'b0;
    assign data[1481] = 16'b0;
    assign data[1482] = ~16'b0;
    assign data[1483] = ~16'b0;
    assign data[1484] = ~16'b0;
    assign data[1485] = ~16'b0;
    assign data[1486] = ~16'b0;
    assign data[1487] = ~16'b0;
    assign data[1488] = ~16'b0;
    assign data[1489] = ~16'b0;
    assign data[1490] = 16'b0;
    assign data[1491] = 16'b0;
    assign data[1492] = ~16'b0;
    assign data[1493] = ~16'b0;
    assign data[1494] = ~16'b0;
    assign data[1495] = ~16'b0;
    assign data[1496] = ~16'b0;
    assign data[1497] = ~16'b0;
    assign data[1498] = ~16'b0;
    assign data[1499] = ~16'b0;
    assign data[1500] = 16'b0;
    assign data[1501] = 16'b0;
    assign data[1502] = ~16'b0;
    assign data[1503] = ~16'b0;
    assign data[1504] = ~16'b0;
    assign data[1505] = ~16'b0;
    assign data[1506] = ~16'b0;
    assign data[1507] = ~16'b0;
    assign data[1508] = ~16'b0;
    assign data[1509] = ~16'b0;
    assign data[1510] = 16'b0;
    assign data[1511] = 16'b0;
    assign data[1512] = ~16'b0;
    assign data[1513] = ~16'b0;
    assign data[1514] = ~16'b0;
    assign data[1515] = ~16'b0;
    assign data[1516] = ~16'b0;
    assign data[1517] = ~16'b0;
    assign data[1518] = ~16'b0;
    assign data[1519] = ~16'b0;
    assign data[1520] = 16'b0;
    assign data[1521] = 16'b0;
    assign data[1522] = ~16'b0;
    assign data[1523] = ~16'b0;
    assign data[1524] = ~16'b0;
    assign data[1525] = ~16'b0;
    assign data[1526] = ~16'b0;
    assign data[1527] = ~16'b0;
    assign data[1528] = ~16'b0;
    assign data[1529] = ~16'b0;
    assign data[1530] = 16'b0;
    assign data[1531] = 16'b0;
    assign data[1532] = ~16'b0;
    assign data[1533] = ~16'b0;
    assign data[1534] = ~16'b0;
    assign data[1535] = ~16'b0;
    assign data[1536] = ~16'b0;
    assign data[1537] = ~16'b0;
    assign data[1538] = ~16'b0;
    assign data[1539] = ~16'b0;
    assign data[1540] = 16'b0;
    assign data[1541] = 16'b0;
    assign data[1542] = ~16'b0;
    assign data[1543] = ~16'b0;
    assign data[1544] = ~16'b0;
    assign data[1545] = ~16'b0;
    assign data[1546] = ~16'b0;
    assign data[1547] = ~16'b0;
    assign data[1548] = ~16'b0;
    assign data[1549] = ~16'b0;
    assign data[1550] = 16'b0;
    assign data[1551] = 16'b0;
    assign data[1552] = ~16'b0;
    assign data[1553] = ~16'b0;
    assign data[1554] = ~16'b0;
    assign data[1555] = ~16'b0;
    assign data[1556] = ~16'b0;
    assign data[1557] = ~16'b0;
    assign data[1558] = ~16'b0;
    assign data[1559] = ~16'b0;
    assign data[1560] = 16'b0;
    assign data[1561] = 16'b0;
    assign data[1562] = ~16'b0;
    assign data[1563] = ~16'b0;
    assign data[1564] = ~16'b0;
    assign data[1565] = ~16'b0;
    assign data[1566] = ~16'b0;
    assign data[1567] = ~16'b0;
    assign data[1568] = ~16'b0;
    assign data[1569] = ~16'b0;
    assign data[1570] = 16'b0;
    assign data[1571] = 16'b0;
    assign data[1572] = ~16'b0;
    assign data[1573] = ~16'b0;
    assign data[1574] = ~16'b0;
    assign data[1575] = ~16'b0;
    assign data[1576] = ~16'b0;
    assign data[1577] = ~16'b0;
    assign data[1578] = ~16'b0;
    assign data[1579] = ~16'b0;
    assign data[1580] = 16'b0;
    assign data[1581] = 16'b0;
    assign data[1582] = ~16'b0;
    assign data[1583] = ~16'b0;
    assign data[1584] = ~16'b0;
    assign data[1585] = ~16'b0;
    assign data[1586] = ~16'b0;
    assign data[1587] = ~16'b0;
    assign data[1588] = ~16'b0;
    assign data[1589] = ~16'b0;
    assign data[1590] = 16'b0;
    assign data[1591] = 16'b0;
    assign data[1592] = ~16'b0;
    assign data[1593] = ~16'b0;
    assign data[1594] = ~16'b0;
    assign data[1595] = ~16'b0;
    assign data[1596] = ~16'b0;
    assign data[1597] = ~16'b0;
    assign data[1598] = ~16'b0;
    assign data[1599] = ~16'b0;
    assign data[1600] = 16'b0;
    assign data[1601] = 16'b0;
    assign data[1602] = ~16'b0;
    assign data[1603] = ~16'b0;
    assign data[1604] = ~16'b0;
    assign data[1605] = ~16'b0;
    assign data[1606] = ~16'b0;
    assign data[1607] = ~16'b0;
    assign data[1608] = ~16'b0;
    assign data[1609] = ~16'b0;
    assign data[1610] = 16'b0;
    assign data[1611] = 16'b0;
    assign data[1612] = ~16'b0;
    assign data[1613] = ~16'b0;
    assign data[1614] = ~16'b0;
    assign data[1615] = ~16'b0;
    assign data[1616] = ~16'b0;
    assign data[1617] = ~16'b0;
    assign data[1618] = ~16'b0;
    assign data[1619] = ~16'b0;
    assign data[1620] = 16'b0;
    assign data[1621] = 16'b0;
    assign data[1622] = ~16'b0;
    assign data[1623] = ~16'b0;
    assign data[1624] = ~16'b0;
    assign data[1625] = ~16'b0;
    assign data[1626] = ~16'b0;
    assign data[1627] = ~16'b0;
    assign data[1628] = ~16'b0;
    assign data[1629] = ~16'b0;
    assign data[1630] = 16'b0;
    assign data[1631] = 16'b0;
    assign data[1632] = ~16'b0;
    assign data[1633] = ~16'b0;
    assign data[1634] = ~16'b0;
    assign data[1635] = ~16'b0;
    assign data[1636] = ~16'b0;
    assign data[1637] = ~16'b0;
    assign data[1638] = ~16'b0;
    assign data[1639] = ~16'b0;
    assign data[1640] = 16'b0;
    assign data[1641] = 16'b0;
    assign data[1642] = ~16'b0;
    assign data[1643] = ~16'b0;
    assign data[1644] = ~16'b0;
    assign data[1645] = ~16'b0;
    assign data[1646] = ~16'b0;
    assign data[1647] = ~16'b0;
    assign data[1648] = ~16'b0;
    assign data[1649] = ~16'b0;
    assign data[1650] = 16'b0;
    assign data[1651] = 16'b0;
    assign data[1652] = ~16'b0;
    assign data[1653] = ~16'b0;
    assign data[1654] = ~16'b0;
    assign data[1655] = ~16'b0;
    assign data[1656] = ~16'b0;
    assign data[1657] = ~16'b0;
    assign data[1658] = ~16'b0;
    assign data[1659] = ~16'b0;
    assign data[1660] = 16'b0;
    assign data[1661] = 16'b0;
    assign data[1662] = ~16'b0;
    assign data[1663] = ~16'b0;
    assign data[1664] = ~16'b0;
    assign data[1665] = ~16'b0;
    assign data[1666] = ~16'b0;
    assign data[1667] = ~16'b0;
    assign data[1668] = ~16'b0;
    assign data[1669] = ~16'b0;
    assign data[1670] = 16'b0;
    assign data[1671] = 16'b0;
    assign data[1672] = ~16'b0;
    assign data[1673] = ~16'b0;
    assign data[1674] = ~16'b0;
    assign data[1675] = ~16'b0;
    assign data[1676] = ~16'b0;
    assign data[1677] = ~16'b0;
    assign data[1678] = ~16'b0;
    assign data[1679] = ~16'b0;
    assign data[1680] = 16'b0;
    assign data[1681] = 16'b0;
    assign data[1682] = ~16'b0;
    assign data[1683] = ~16'b0;
    assign data[1684] = ~16'b0;
    assign data[1685] = ~16'b0;
    assign data[1686] = ~16'b0;
    assign data[1687] = ~16'b0;
    assign data[1688] = ~16'b0;
    assign data[1689] = ~16'b0;
    assign data[1690] = 16'b0;
    assign data[1691] = 16'b0;
    assign data[1692] = ~16'b0;
    assign data[1693] = ~16'b0;
    assign data[1694] = ~16'b0;
    assign data[1695] = ~16'b0;
    assign data[1696] = ~16'b0;
    assign data[1697] = ~16'b0;
    assign data[1698] = ~16'b0;
    assign data[1699] = ~16'b0;
    assign data[1700] = 16'b0;
    assign data[1701] = 16'b0;
    assign data[1702] = ~16'b0;
    assign data[1703] = ~16'b0;
    assign data[1704] = ~16'b0;
    assign data[1705] = ~16'b0;
    assign data[1706] = ~16'b0;
    assign data[1707] = ~16'b0;
    assign data[1708] = ~16'b0;
    assign data[1709] = ~16'b0;
    assign data[1710] = 16'b0;
    assign data[1711] = 16'b0;
    assign data[1712] = ~16'b0;
    assign data[1713] = ~16'b0;
    assign data[1714] = ~16'b0;
    assign data[1715] = ~16'b0;
    assign data[1716] = ~16'b0;
    assign data[1717] = ~16'b0;
    assign data[1718] = ~16'b0;
    assign data[1719] = ~16'b0;
    assign data[1720] = 16'b0;
    assign data[1721] = 16'b0;
    assign data[1722] = ~16'b0;
    assign data[1723] = ~16'b0;
    assign data[1724] = ~16'b0;
    assign data[1725] = ~16'b0;
    assign data[1726] = ~16'b0;
    assign data[1727] = ~16'b0;
    assign data[1728] = ~16'b0;
    assign data[1729] = ~16'b0;
    assign data[1730] = 16'b0;
    assign data[1731] = 16'b0;
    assign data[1732] = ~16'b0;
    assign data[1733] = ~16'b0;
    assign data[1734] = ~16'b0;
    assign data[1735] = ~16'b0;
    assign data[1736] = ~16'b0;
    assign data[1737] = ~16'b0;
    assign data[1738] = ~16'b0;
    assign data[1739] = ~16'b0;
    assign data[1740] = 16'b0;
    assign data[1741] = 16'b0;
    assign data[1742] = ~16'b0;
    assign data[1743] = ~16'b0;
    assign data[1744] = ~16'b0;
    assign data[1745] = ~16'b0;
    assign data[1746] = ~16'b0;
    assign data[1747] = ~16'b0;
    assign data[1748] = ~16'b0;
    assign data[1749] = ~16'b0;
    assign data[1750] = 16'b0;
    assign data[1751] = 16'b0;
    assign data[1752] = ~16'b0;
    assign data[1753] = ~16'b0;
    assign data[1754] = ~16'b0;
    assign data[1755] = ~16'b0;
    assign data[1756] = ~16'b0;
    assign data[1757] = ~16'b0;
    assign data[1758] = ~16'b0;
    assign data[1759] = ~16'b0;
    assign data[1760] = 16'b0;
    assign data[1761] = 16'b0;
    assign data[1762] = ~16'b0;
    assign data[1763] = ~16'b0;
    assign data[1764] = ~16'b0;
    assign data[1765] = ~16'b0;
    assign data[1766] = ~16'b0;
    assign data[1767] = ~16'b0;
    assign data[1768] = ~16'b0;
    assign data[1769] = ~16'b0;
    assign data[1770] = 16'b0;
    assign data[1771] = 16'b0;
    assign data[1772] = ~16'b0;
    assign data[1773] = ~16'b0;
    assign data[1774] = ~16'b0;
    assign data[1775] = ~16'b0;
    assign data[1776] = ~16'b0;
    assign data[1777] = ~16'b0;
    assign data[1778] = ~16'b0;
    assign data[1779] = ~16'b0;
    assign data[1780] = 16'b0;
    assign data[1781] = 16'b0;
    assign data[1782] = ~16'b0;
    assign data[1783] = ~16'b0;
    assign data[1784] = ~16'b0;
    assign data[1785] = ~16'b0;
    assign data[1786] = ~16'b0;
    assign data[1787] = ~16'b0;
    assign data[1788] = ~16'b0;
    assign data[1789] = ~16'b0;
    assign data[1790] = 16'b0;
    assign data[1791] = 16'b0;
    assign data[1792] = ~16'b0;
    assign data[1793] = ~16'b0;
    assign data[1794] = ~16'b0;
    assign data[1795] = ~16'b0;
    assign data[1796] = ~16'b0;
    assign data[1797] = ~16'b0;
    assign data[1798] = ~16'b0;
    assign data[1799] = ~16'b0;
    assign data[1800] = 16'b0;
    assign data[1801] = 16'b0;
    assign data[1802] = ~16'b0;
    assign data[1803] = ~16'b0;
    assign data[1804] = ~16'b0;
    assign data[1805] = ~16'b0;
    assign data[1806] = ~16'b0;
    assign data[1807] = ~16'b0;
    assign data[1808] = ~16'b0;
    assign data[1809] = ~16'b0;
    assign data[1810] = 16'b0;
    assign data[1811] = 16'b0;
    assign data[1812] = ~16'b0;
    assign data[1813] = ~16'b0;
    assign data[1814] = ~16'b0;
    assign data[1815] = ~16'b0;
    assign data[1816] = ~16'b0;
    assign data[1817] = ~16'b0;
    assign data[1818] = ~16'b0;
    assign data[1819] = ~16'b0;
    assign data[1820] = 16'b0;
    assign data[1821] = 16'b0;
    assign data[1822] = ~16'b0;
    assign data[1823] = ~16'b0;
    assign data[1824] = ~16'b0;
    assign data[1825] = ~16'b0;
    assign data[1826] = ~16'b0;
    assign data[1827] = ~16'b0;
    assign data[1828] = ~16'b0;
    assign data[1829] = ~16'b0;
    assign data[1830] = 16'b0;
    assign data[1831] = 16'b0;
    assign data[1832] = ~16'b0;
    assign data[1833] = ~16'b0;
    assign data[1834] = ~16'b0;
    assign data[1835] = ~16'b0;
    assign data[1836] = ~16'b0;
    assign data[1837] = ~16'b0;
    assign data[1838] = ~16'b0;
    assign data[1839] = ~16'b0;
    assign data[1840] = 16'b0;
    assign data[1841] = 16'b0;
    assign data[1842] = ~16'b0;
    assign data[1843] = ~16'b0;
    assign data[1844] = ~16'b0;
    assign data[1845] = ~16'b0;
    assign data[1846] = ~16'b0;
    assign data[1847] = ~16'b0;
    assign data[1848] = ~16'b0;
    assign data[1849] = ~16'b0;
    assign data[1850] = 16'b0;
    assign data[1851] = 16'b0;
    assign data[1852] = ~16'b0;
    assign data[1853] = ~16'b0;
    assign data[1854] = ~16'b0;
    assign data[1855] = ~16'b0;
    assign data[1856] = ~16'b0;
    assign data[1857] = ~16'b0;
    assign data[1858] = ~16'b0;
    assign data[1859] = ~16'b0;
    assign data[1860] = 16'b0;
    assign data[1861] = 16'b0;
    assign data[1862] = ~16'b0;
    assign data[1863] = ~16'b0;
    assign data[1864] = ~16'b0;
    assign data[1865] = ~16'b0;
    assign data[1866] = ~16'b0;
    assign data[1867] = ~16'b0;
    assign data[1868] = ~16'b0;
    assign data[1869] = ~16'b0;
    assign data[1870] = 16'b0;
    assign data[1871] = 16'b0;
    assign data[1872] = 16'b0;
    assign data[1873] = 16'b0;
    assign data[1874] = 16'b0;
    assign data[1875] = 16'b0;
    assign data[1876] = 16'b0;
    assign data[1877] = 16'b0;
    assign data[1878] = 16'b0;
    assign data[1879] = 16'b0;
    assign data[1880] = 16'b0;
    assign data[1881] = 16'b0;
    assign data[1882] = 16'b0;
    assign data[1883] = 16'b0;
    assign data[1884] = 16'b0;
    assign data[1885] = 16'b0;
    assign data[1886] = 16'b0;
    assign data[1887] = 16'b0;
    assign data[1888] = 16'b0;
    assign data[1889] = 16'b0;
    assign data[1890] = ~16'b0;
    assign data[1891] = ~16'b0;
    assign data[1892] = ~16'b0;
    assign data[1893] = ~16'b0;
    assign data[1894] = ~16'b0;
    assign data[1895] = ~16'b0;
    assign data[1896] = ~16'b0;
    assign data[1897] = ~16'b0;
    assign data[1898] = ~16'b0;
    assign data[1899] = ~16'b0;
    assign data[1900] = ~16'b0;
    assign data[1901] = ~16'b0;
    assign data[1902] = ~16'b0;
    assign data[1903] = ~16'b0;
    assign data[1904] = ~16'b0;
    assign data[1905] = ~16'b0;
    assign data[1906] = ~16'b0;
    assign data[1907] = ~16'b0;
    assign data[1908] = ~16'b0;
    assign data[1909] = ~16'b0;
    assign data[1910] = ~16'b0;
    assign data[1911] = ~16'b0;
    assign data[1912] = ~16'b0;
    assign data[1913] = ~16'b0;
    assign data[1914] = ~16'b0;
    assign data[1915] = ~16'b0;
    assign data[1916] = ~16'b0;
    assign data[1917] = ~16'b0;
    assign data[1918] = ~16'b0;
    assign data[1919] = ~16'b0;
    assign data[1920] = ~16'b0;
    assign data[1921] = ~16'b0;
    assign data[1922] = ~16'b0;
    assign data[1923] = ~16'b0;
    assign data[1924] = ~16'b0;
    assign data[1925] = ~16'b0;
    assign data[1926] = ~16'b0;
    assign data[1927] = ~16'b0;
    assign data[1928] = ~16'b0;
    assign data[1929] = ~16'b0;
    assign data[1930] = ~16'b0;
    assign data[1931] = ~16'b0;
    assign data[1932] = ~16'b0;
    assign data[1933] = ~16'b0;
    assign data[1934] = ~16'b0;
    assign data[1935] = ~16'b0;
    assign data[1936] = ~16'b0;
    assign data[1937] = ~16'b0;
    assign data[1938] = ~16'b0;
    assign data[1939] = ~16'b0;
    assign data[1940] = ~16'b0;
    assign data[1941] = ~16'b0;
    assign data[1942] = ~16'b0;
    assign data[1943] = ~16'b0;
    assign data[1944] = ~16'b0;
    assign data[1945] = ~16'b0;
    assign data[1946] = ~16'b0;
    assign data[1947] = ~16'b0;
    assign data[1948] = ~16'b0;
    assign data[1949] = ~16'b0;
    assign data[1950] = ~16'b0;
    assign data[1951] = ~16'b0;
    assign data[1952] = ~16'b0;
    assign data[1953] = ~16'b0;
    assign data[1954] = ~16'b0;
    assign data[1955] = ~16'b0;
    assign data[1956] = ~16'b0;
    assign data[1957] = ~16'b0;
    assign data[1958] = ~16'b0;
    assign data[1959] = ~16'b0;
    assign data[1960] = ~16'b0;
    assign data[1961] = ~16'b0;
    assign data[1962] = ~16'b0;
    assign data[1963] = ~16'b0;
    assign data[1964] = ~16'b0;
    assign data[1965] = ~16'b0;
    assign data[1966] = ~16'b0;
    assign data[1967] = ~16'b0;
    assign data[1968] = ~16'b0;
    assign data[1969] = ~16'b0;
    assign data[1970] = ~16'b0;
    assign data[1971] = ~16'b0;
    assign data[1972] = ~16'b0;
    assign data[1973] = ~16'b0;
    assign data[1974] = ~16'b0;
    assign data[1975] = ~16'b0;
    assign data[1976] = ~16'b0;
    assign data[1977] = ~16'b0;
    assign data[1978] = ~16'b0;
    assign data[1979] = ~16'b0;
    assign data[1980] = ~16'b0;
    assign data[1981] = ~16'b0;
    assign data[1982] = ~16'b0;
    assign data[1983] = ~16'b0;
    assign data[1984] = ~16'b0;
    assign data[1985] = ~16'b0;
    assign data[1986] = ~16'b0;
    assign data[1987] = ~16'b0;
    assign data[1988] = ~16'b0;
    assign data[1989] = ~16'b0;
    assign data[1990] = ~16'b0;
    assign data[1991] = ~16'b0;
    assign data[1992] = ~16'b0;
    assign data[1993] = ~16'b0;
    assign data[1994] = ~16'b0;
    assign data[1995] = ~16'b0;
    assign data[1996] = ~16'b0;
    assign data[1997] = ~16'b0;
    assign data[1998] = ~16'b0;
    assign data[1999] = ~16'b0;
    assign data[2000] = ~16'b0;
    assign data[2001] = ~16'b0;
    assign data[2002] = ~16'b0;
    assign data[2003] = ~16'b0;
    assign data[2004] = ~16'b0;
    assign data[2005] = ~16'b0;
    assign data[2006] = ~16'b0;
    assign data[2007] = ~16'b0;
    assign data[2008] = ~16'b0;
    assign data[2009] = ~16'b0;
    assign data[2010] = ~16'b0;
    assign data[2011] = ~16'b0;
    assign data[2012] = ~16'b0;
    assign data[2013] = ~16'b0;
    assign data[2014] = ~16'b0;
    assign data[2015] = ~16'b0;
    assign data[2016] = ~16'b0;
    assign data[2017] = ~16'b0;
    assign data[2018] = ~16'b0;
    assign data[2019] = ~16'b0;
    assign data[2020] = ~16'b0;
    assign data[2021] = ~16'b0;
    assign data[2022] = ~16'b0;
    assign data[2023] = ~16'b0;
    assign data[2024] = ~16'b0;
    assign data[2025] = ~16'b0;
    assign data[2026] = ~16'b0;
    assign data[2027] = ~16'b0;
    assign data[2028] = ~16'b0;
    assign data[2029] = ~16'b0;
    assign data[2030] = ~16'b0;
    assign data[2031] = ~16'b0;
    assign data[2032] = ~16'b0;
    assign data[2033] = ~16'b0;
    assign data[2034] = ~16'b0;
    assign data[2035] = ~16'b0;
    assign data[2036] = ~16'b0;
    assign data[2037] = ~16'b0;
    assign data[2038] = ~16'b0;
    assign data[2039] = ~16'b0;
    assign data[2040] = ~16'b0;
    assign data[2041] = ~16'b0;
    assign data[2042] = ~16'b0;
    assign data[2043] = ~16'b0;
    assign data[2044] = ~16'b0;
    assign data[2045] = ~16'b0;
    assign data[2046] = ~16'b0;
    assign data[2047] = ~16'b0;
    assign data[2048] = ~16'b0;
    assign data[2049] = ~16'b0;
    assign data[2050] = ~16'b0;
    assign data[2051] = ~16'b0;
    assign data[2052] = ~16'b0;
    assign data[2053] = ~16'b0;
    assign data[2054] = ~16'b0;
    assign data[2055] = ~16'b0;
    assign data[2056] = ~16'b0;
    assign data[2057] = ~16'b0;
    assign data[2058] = ~16'b0;
    assign data[2059] = ~16'b0;
    assign data[2060] = ~16'b0;
    assign data[2061] = ~16'b0;
    assign data[2062] = ~16'b0;
    assign data[2063] = ~16'b0;
    assign data[2064] = ~16'b0;
    assign data[2065] = ~16'b0;
    assign data[2066] = ~16'b0;
    assign data[2067] = ~16'b0;
    assign data[2068] = ~16'b0;
    assign data[2069] = ~16'b0;
    assign data[2070] = 16'b0;
    assign data[2071] = 16'b0;
    assign data[2072] = 16'b0;
    assign data[2073] = 16'b0;
    assign data[2074] = 16'b0;
    assign data[2075] = 16'b0;
    assign data[2076] = 16'b0;
    assign data[2077] = 16'b0;
    assign data[2078] = 16'b0;
    assign data[2079] = 16'b0;
    assign data[2080] = 16'b0;
    assign data[2081] = 16'b0;
    assign data[2082] = 16'b0;
    assign data[2083] = 16'b0;
    assign data[2084] = 16'b0;
    assign data[2085] = 16'b0;
    assign data[2086] = 16'b0;
    assign data[2087] = 16'b0;
    assign data[2088] = 16'b0;
    assign data[2089] = 16'b0;
    assign data[2090] = 16'b0;
    assign data[2091] = 16'b0;
    assign data[2092] = ~16'b0;
    assign data[2093] = ~16'b0;
    assign data[2094] = ~16'b0;
    assign data[2095] = ~16'b0;
    assign data[2096] = ~16'b0;
    assign data[2097] = ~16'b0;
    assign data[2098] = ~16'b0;
    assign data[2099] = ~16'b0;
    assign data[2100] = 16'b0;
    assign data[2101] = 16'b0;
    assign data[2102] = ~16'b0;
    assign data[2103] = ~16'b0;
    assign data[2104] = ~16'b0;
    assign data[2105] = ~16'b0;
    assign data[2106] = ~16'b0;
    assign data[2107] = ~16'b0;
    assign data[2108] = ~16'b0;
    assign data[2109] = ~16'b0;
    assign data[2110] = 16'b0;
    assign data[2111] = 16'b0;
    assign data[2112] = ~16'b0;
    assign data[2113] = ~16'b0;
    assign data[2114] = ~16'b0;
    assign data[2115] = ~16'b0;
    assign data[2116] = ~16'b0;
    assign data[2117] = ~16'b0;
    assign data[2118] = ~16'b0;
    assign data[2119] = ~16'b0;
    assign data[2120] = 16'b0;
    assign data[2121] = 16'b0;
    assign data[2122] = ~16'b0;
    assign data[2123] = ~16'b0;
    assign data[2124] = ~16'b0;
    assign data[2125] = ~16'b0;
    assign data[2126] = ~16'b0;
    assign data[2127] = ~16'b0;
    assign data[2128] = ~16'b0;
    assign data[2129] = ~16'b0;
    assign data[2130] = 16'b0;
    assign data[2131] = 16'b0;
    assign data[2132] = ~16'b0;
    assign data[2133] = ~16'b0;
    assign data[2134] = ~16'b0;
    assign data[2135] = ~16'b0;
    assign data[2136] = ~16'b0;
    assign data[2137] = ~16'b0;
    assign data[2138] = ~16'b0;
    assign data[2139] = ~16'b0;
    assign data[2140] = 16'b0;
    assign data[2141] = 16'b0;
    assign data[2142] = ~16'b0;
    assign data[2143] = ~16'b0;
    assign data[2144] = ~16'b0;
    assign data[2145] = ~16'b0;
    assign data[2146] = ~16'b0;
    assign data[2147] = ~16'b0;
    assign data[2148] = ~16'b0;
    assign data[2149] = ~16'b0;
    assign data[2150] = 16'b0;
    assign data[2151] = 16'b0;
    assign data[2152] = ~16'b0;
    assign data[2153] = ~16'b0;
    assign data[2154] = ~16'b0;
    assign data[2155] = ~16'b0;
    assign data[2156] = ~16'b0;
    assign data[2157] = ~16'b0;
    assign data[2158] = ~16'b0;
    assign data[2159] = ~16'b0;
    assign data[2160] = 16'b0;
    assign data[2161] = 16'b0;
    assign data[2162] = ~16'b0;
    assign data[2163] = ~16'b0;
    assign data[2164] = ~16'b0;
    assign data[2165] = ~16'b0;
    assign data[2166] = ~16'b0;
    assign data[2167] = ~16'b0;
    assign data[2168] = ~16'b0;
    assign data[2169] = ~16'b0;
    assign data[2170] = 16'b0;
    assign data[2171] = 16'b0;
    assign data[2172] = ~16'b0;
    assign data[2173] = ~16'b0;
    assign data[2174] = ~16'b0;
    assign data[2175] = ~16'b0;
    assign data[2176] = ~16'b0;
    assign data[2177] = ~16'b0;
    assign data[2178] = ~16'b0;
    assign data[2179] = ~16'b0;
    assign data[2180] = 16'b0;
    assign data[2181] = 16'b0;
    assign data[2182] = ~16'b0;
    assign data[2183] = ~16'b0;
    assign data[2184] = ~16'b0;
    assign data[2185] = ~16'b0;
    assign data[2186] = ~16'b0;
    assign data[2187] = ~16'b0;
    assign data[2188] = ~16'b0;
    assign data[2189] = ~16'b0;
    assign data[2190] = 16'b0;
    assign data[2191] = 16'b0;
    assign data[2192] = ~16'b0;
    assign data[2193] = ~16'b0;
    assign data[2194] = ~16'b0;
    assign data[2195] = ~16'b0;
    assign data[2196] = ~16'b0;
    assign data[2197] = ~16'b0;
    assign data[2198] = ~16'b0;
    assign data[2199] = ~16'b0;
    assign data[2200] = 16'b0;
    assign data[2201] = 16'b0;
    assign data[2202] = ~16'b0;
    assign data[2203] = ~16'b0;
    assign data[2204] = ~16'b0;
    assign data[2205] = ~16'b0;
    assign data[2206] = ~16'b0;
    assign data[2207] = ~16'b0;
    assign data[2208] = ~16'b0;
    assign data[2209] = ~16'b0;
    assign data[2210] = 16'b0;
    assign data[2211] = 16'b0;
    assign data[2212] = ~16'b0;
    assign data[2213] = ~16'b0;
    assign data[2214] = ~16'b0;
    assign data[2215] = ~16'b0;
    assign data[2216] = ~16'b0;
    assign data[2217] = ~16'b0;
    assign data[2218] = ~16'b0;
    assign data[2219] = ~16'b0;
    assign data[2220] = 16'b0;
    assign data[2221] = 16'b0;
    assign data[2222] = ~16'b0;
    assign data[2223] = ~16'b0;
    assign data[2224] = ~16'b0;
    assign data[2225] = ~16'b0;
    assign data[2226] = ~16'b0;
    assign data[2227] = ~16'b0;
    assign data[2228] = ~16'b0;
    assign data[2229] = ~16'b0;
    assign data[2230] = 16'b0;
    assign data[2231] = 16'b0;
    assign data[2232] = ~16'b0;
    assign data[2233] = ~16'b0;
    assign data[2234] = ~16'b0;
    assign data[2235] = ~16'b0;
    assign data[2236] = ~16'b0;
    assign data[2237] = ~16'b0;
    assign data[2238] = ~16'b0;
    assign data[2239] = ~16'b0;
    assign data[2240] = 16'b0;
    assign data[2241] = 16'b0;
    assign data[2242] = ~16'b0;
    assign data[2243] = ~16'b0;
    assign data[2244] = ~16'b0;
    assign data[2245] = ~16'b0;
    assign data[2246] = ~16'b0;
    assign data[2247] = ~16'b0;
    assign data[2248] = ~16'b0;
    assign data[2249] = ~16'b0;
    assign data[2250] = 16'b0;
    assign data[2251] = 16'b0;
    assign data[2252] = ~16'b0;
    assign data[2253] = ~16'b0;
    assign data[2254] = ~16'b0;
    assign data[2255] = ~16'b0;
    assign data[2256] = ~16'b0;
    assign data[2257] = ~16'b0;
    assign data[2258] = ~16'b0;
    assign data[2259] = ~16'b0;
    assign data[2260] = 16'b0;
    assign data[2261] = 16'b0;
    assign data[2262] = ~16'b0;
    assign data[2263] = ~16'b0;
    assign data[2264] = ~16'b0;
    assign data[2265] = ~16'b0;
    assign data[2266] = ~16'b0;
    assign data[2267] = ~16'b0;
    assign data[2268] = ~16'b0;
    assign data[2269] = ~16'b0;
    assign data[2270] = 16'b0;
    assign data[2271] = 16'b0;
    assign data[2272] = ~16'b0;
    assign data[2273] = ~16'b0;
    assign data[2274] = ~16'b0;
    assign data[2275] = ~16'b0;
    assign data[2276] = ~16'b0;
    assign data[2277] = ~16'b0;
    assign data[2278] = ~16'b0;
    assign data[2279] = ~16'b0;
    assign data[2280] = 16'b0;
    assign data[2281] = 16'b0;
    assign data[2282] = ~16'b0;
    assign data[2283] = ~16'b0;
    assign data[2284] = ~16'b0;
    assign data[2285] = ~16'b0;
    assign data[2286] = ~16'b0;
    assign data[2287] = ~16'b0;
    assign data[2288] = ~16'b0;
    assign data[2289] = ~16'b0;
    assign data[2290] = 16'b0;
    assign data[2291] = 16'b0;
    assign data[2292] = ~16'b0;
    assign data[2293] = ~16'b0;
    assign data[2294] = ~16'b0;
    assign data[2295] = ~16'b0;
    assign data[2296] = ~16'b0;
    assign data[2297] = ~16'b0;
    assign data[2298] = ~16'b0;
    assign data[2299] = ~16'b0;
    assign data[2300] = 16'b0;
    assign data[2301] = 16'b0;
    assign data[2302] = ~16'b0;
    assign data[2303] = ~16'b0;
    assign data[2304] = ~16'b0;
    assign data[2305] = ~16'b0;
    assign data[2306] = ~16'b0;
    assign data[2307] = ~16'b0;
    assign data[2308] = ~16'b0;
    assign data[2309] = ~16'b0;
    assign data[2310] = 16'b0;
    assign data[2311] = 16'b0;
    assign data[2312] = ~16'b0;
    assign data[2313] = ~16'b0;
    assign data[2314] = ~16'b0;
    assign data[2315] = ~16'b0;
    assign data[2316] = ~16'b0;
    assign data[2317] = ~16'b0;
    assign data[2318] = ~16'b0;
    assign data[2319] = ~16'b0;
    assign data[2320] = 16'b0;
    assign data[2321] = 16'b0;
    assign data[2322] = ~16'b0;
    assign data[2323] = ~16'b0;
    assign data[2324] = ~16'b0;
    assign data[2325] = ~16'b0;
    assign data[2326] = ~16'b0;
    assign data[2327] = ~16'b0;
    assign data[2328] = ~16'b0;
    assign data[2329] = ~16'b0;
    assign data[2330] = 16'b0;
    assign data[2331] = 16'b0;
    assign data[2332] = ~16'b0;
    assign data[2333] = ~16'b0;
    assign data[2334] = ~16'b0;
    assign data[2335] = ~16'b0;
    assign data[2336] = ~16'b0;
    assign data[2337] = ~16'b0;
    assign data[2338] = ~16'b0;
    assign data[2339] = ~16'b0;
    assign data[2340] = 16'b0;
    assign data[2341] = 16'b0;
    assign data[2342] = ~16'b0;
    assign data[2343] = ~16'b0;
    assign data[2344] = ~16'b0;
    assign data[2345] = ~16'b0;
    assign data[2346] = ~16'b0;
    assign data[2347] = ~16'b0;
    assign data[2348] = ~16'b0;
    assign data[2349] = ~16'b0;
    assign data[2350] = 16'b0;
    assign data[2351] = 16'b0;
    assign data[2352] = ~16'b0;
    assign data[2353] = ~16'b0;
    assign data[2354] = ~16'b0;
    assign data[2355] = ~16'b0;
    assign data[2356] = ~16'b0;
    assign data[2357] = ~16'b0;
    assign data[2358] = ~16'b0;
    assign data[2359] = ~16'b0;
    assign data[2360] = 16'b0;
    assign data[2361] = 16'b0;
    assign data[2362] = ~16'b0;
    assign data[2363] = ~16'b0;
    assign data[2364] = ~16'b0;
    assign data[2365] = ~16'b0;
    assign data[2366] = ~16'b0;
    assign data[2367] = ~16'b0;
    assign data[2368] = ~16'b0;
    assign data[2369] = ~16'b0;
    assign data[2370] = 16'b0;
    assign data[2371] = 16'b0;
    assign data[2372] = ~16'b0;
    assign data[2373] = ~16'b0;
    assign data[2374] = ~16'b0;
    assign data[2375] = ~16'b0;
    assign data[2376] = ~16'b0;
    assign data[2377] = ~16'b0;
    assign data[2378] = ~16'b0;
    assign data[2379] = ~16'b0;
    assign data[2380] = 16'b0;
    assign data[2381] = 16'b0;
    assign data[2382] = ~16'b0;
    assign data[2383] = ~16'b0;
    assign data[2384] = ~16'b0;
    assign data[2385] = ~16'b0;
    assign data[2386] = ~16'b0;
    assign data[2387] = ~16'b0;
    assign data[2388] = ~16'b0;
    assign data[2389] = ~16'b0;
    assign data[2390] = 16'b0;
    assign data[2391] = 16'b0;
    assign data[2392] = ~16'b0;
    assign data[2393] = ~16'b0;
    assign data[2394] = ~16'b0;
    assign data[2395] = ~16'b0;
    assign data[2396] = ~16'b0;
    assign data[2397] = ~16'b0;
    assign data[2398] = ~16'b0;
    assign data[2399] = ~16'b0;
    assign data[2400] = 16'b0;
    assign data[2401] = 16'b0;
    assign data[2402] = ~16'b0;
    assign data[2403] = ~16'b0;
    assign data[2404] = ~16'b0;
    assign data[2405] = ~16'b0;
    assign data[2406] = ~16'b0;
    assign data[2407] = ~16'b0;
    assign data[2408] = ~16'b0;
    assign data[2409] = ~16'b0;
    assign data[2410] = 16'b0;
    assign data[2411] = 16'b0;
    assign data[2412] = ~16'b0;
    assign data[2413] = ~16'b0;
    assign data[2414] = ~16'b0;
    assign data[2415] = ~16'b0;
    assign data[2416] = ~16'b0;
    assign data[2417] = ~16'b0;
    assign data[2418] = ~16'b0;
    assign data[2419] = ~16'b0;
    assign data[2420] = 16'b0;
    assign data[2421] = 16'b0;
    assign data[2422] = ~16'b0;
    assign data[2423] = ~16'b0;
    assign data[2424] = ~16'b0;
    assign data[2425] = ~16'b0;
    assign data[2426] = ~16'b0;
    assign data[2427] = ~16'b0;
    assign data[2428] = ~16'b0;
    assign data[2429] = ~16'b0;
    assign data[2430] = 16'b0;
    assign data[2431] = 16'b0;
    assign data[2432] = ~16'b0;
    assign data[2433] = ~16'b0;
    assign data[2434] = ~16'b0;
    assign data[2435] = ~16'b0;
    assign data[2436] = ~16'b0;
    assign data[2437] = ~16'b0;
    assign data[2438] = ~16'b0;
    assign data[2439] = ~16'b0;
    assign data[2440] = 16'b0;
    assign data[2441] = 16'b0;
    assign data[2442] = 16'b0;
    assign data[2443] = 16'b0;
    assign data[2444] = 16'b0;
    assign data[2445] = 16'b0;
    assign data[2446] = 16'b0;
    assign data[2447] = 16'b0;
    assign data[2448] = 16'b0;
    assign data[2449] = 16'b0;
    assign data[2450] = 16'b0;
    assign data[2451] = 16'b0;
    assign data[2452] = 16'b0;
    assign data[2453] = 16'b0;
    assign data[2454] = 16'b0;
    assign data[2455] = 16'b0;
    assign data[2456] = 16'b0;
    assign data[2457] = 16'b0;
    assign data[2458] = 16'b0;
    assign data[2459] = 16'b0;
    assign data[2460] = ~16'b0;
    assign data[2461] = ~16'b0;
    assign data[2462] = ~16'b0;
    assign data[2463] = ~16'b0;
    assign data[2464] = ~16'b0;
    assign data[2465] = ~16'b0;
    assign data[2466] = ~16'b0;
    assign data[2467] = ~16'b0;
    assign data[2468] = ~16'b0;
    assign data[2469] = ~16'b0;
    assign data[2470] = ~16'b0;
    assign data[2471] = ~16'b0;
    assign data[2472] = ~16'b0;
    assign data[2473] = ~16'b0;
    assign data[2474] = ~16'b0;
    assign data[2475] = ~16'b0;
    assign data[2476] = ~16'b0;
    assign data[2477] = ~16'b0;
    assign data[2478] = ~16'b0;
    assign data[2479] = ~16'b0;
    assign data[2480] = ~16'b0;
    assign data[2481] = ~16'b0;
    assign data[2482] = ~16'b0;
    assign data[2483] = ~16'b0;
    assign data[2484] = ~16'b0;
    assign data[2485] = ~16'b0;
    assign data[2486] = ~16'b0;
    assign data[2487] = ~16'b0;
    assign data[2488] = ~16'b0;
    assign data[2489] = ~16'b0;
    assign data[2490] = ~16'b0;
    assign data[2491] = ~16'b0;
    assign data[2492] = ~16'b0;
    assign data[2493] = ~16'b0;
    assign data[2494] = ~16'b0;
    assign data[2495] = ~16'b0;
    assign data[2496] = ~16'b0;
    assign data[2497] = ~16'b0;
    assign data[2498] = ~16'b0;
    assign data[2499] = ~16'b0;
    assign data[2500] = ~16'b0;
    assign data[2501] = ~16'b0;
    assign data[2502] = ~16'b0;
    assign data[2503] = ~16'b0;
    assign data[2504] = ~16'b0;
    assign data[2505] = ~16'b0;
    assign data[2506] = ~16'b0;
    assign data[2507] = ~16'b0;
    assign data[2508] = ~16'b0;
    assign data[2509] = ~16'b0;
    assign data[2510] = ~16'b0;
    assign data[2511] = ~16'b0;
    assign data[2512] = ~16'b0;
    assign data[2513] = ~16'b0;
    assign data[2514] = ~16'b0;
    assign data[2515] = ~16'b0;
    assign data[2516] = ~16'b0;
    assign data[2517] = ~16'b0;
    assign data[2518] = ~16'b0;
    assign data[2519] = ~16'b0;
    assign data[2520] = ~16'b0;
    assign data[2521] = ~16'b0;
    assign data[2522] = ~16'b0;
    assign data[2523] = ~16'b0;
    assign data[2524] = ~16'b0;
    assign data[2525] = ~16'b0;
    assign data[2526] = ~16'b0;
    assign data[2527] = ~16'b0;
    assign data[2528] = ~16'b0;
    assign data[2529] = ~16'b0;
    assign data[2530] = ~16'b0;
    assign data[2531] = ~16'b0;
    assign data[2532] = ~16'b0;
    assign data[2533] = ~16'b0;
    assign data[2534] = ~16'b0;
    assign data[2535] = ~16'b0;
    assign data[2536] = ~16'b0;
    assign data[2537] = ~16'b0;
    assign data[2538] = ~16'b0;
    assign data[2539] = ~16'b0;
    assign data[2540] = ~16'b0;
    assign data[2541] = ~16'b0;
    assign data[2542] = ~16'b0;
    assign data[2543] = ~16'b0;
    assign data[2544] = ~16'b0;
    assign data[2545] = ~16'b0;
    assign data[2546] = ~16'b0;
    assign data[2547] = ~16'b0;
    assign data[2548] = ~16'b0;
    assign data[2549] = ~16'b0;
    assign data[2550] = ~16'b0;
    assign data[2551] = ~16'b0;
    assign data[2552] = ~16'b0;
    assign data[2553] = ~16'b0;
    assign data[2554] = ~16'b0;
    assign data[2555] = ~16'b0;
    assign data[2556] = ~16'b0;
    assign data[2557] = ~16'b0;
    assign data[2558] = ~16'b0;
    assign data[2559] = ~16'b0;
    assign data[2560] = ~16'b0;
    assign data[2561] = ~16'b0;
    assign data[2562] = ~16'b0;
    assign data[2563] = ~16'b0;
    assign data[2564] = ~16'b0;
    assign data[2565] = ~16'b0;
    assign data[2566] = ~16'b0;
    assign data[2567] = ~16'b0;
    assign data[2568] = ~16'b0;
    assign data[2569] = ~16'b0;
    assign data[2570] = ~16'b0;
    assign data[2571] = ~16'b0;
    assign data[2572] = ~16'b0;
    assign data[2573] = ~16'b0;
    assign data[2574] = ~16'b0;
    assign data[2575] = ~16'b0;
    assign data[2576] = ~16'b0;
    assign data[2577] = ~16'b0;
    assign data[2578] = ~16'b0;
    assign data[2579] = ~16'b0;
    assign data[2580] = ~16'b0;
    assign data[2581] = ~16'b0;
    assign data[2582] = ~16'b0;
    assign data[2583] = ~16'b0;
    assign data[2584] = ~16'b0;
    assign data[2585] = ~16'b0;
    assign data[2586] = ~16'b0;
    assign data[2587] = ~16'b0;
    assign data[2588] = ~16'b0;
    assign data[2589] = ~16'b0;
    assign data[2590] = ~16'b0;
    assign data[2591] = ~16'b0;
    assign data[2592] = ~16'b0;
    assign data[2593] = ~16'b0;
    assign data[2594] = ~16'b0;
    assign data[2595] = ~16'b0;
    assign data[2596] = ~16'b0;
    assign data[2597] = ~16'b0;
    assign data[2598] = ~16'b0;
    assign data[2599] = ~16'b0;
    assign data[2600] = ~16'b0;
    assign data[2601] = ~16'b0;
    assign data[2602] = ~16'b0;
    assign data[2603] = ~16'b0;
    assign data[2604] = ~16'b0;
    assign data[2605] = ~16'b0;
    assign data[2606] = ~16'b0;
    assign data[2607] = ~16'b0;
    assign data[2608] = ~16'b0;
    assign data[2609] = ~16'b0;
    assign data[2610] = ~16'b0;
    assign data[2611] = ~16'b0;
    assign data[2612] = ~16'b0;
    assign data[2613] = ~16'b0;
    assign data[2614] = ~16'b0;
    assign data[2615] = ~16'b0;
    assign data[2616] = ~16'b0;
    assign data[2617] = ~16'b0;
    assign data[2618] = ~16'b0;
    assign data[2619] = ~16'b0;
    assign data[2620] = ~16'b0;
    assign data[2621] = ~16'b0;
    assign data[2622] = ~16'b0;
    assign data[2623] = ~16'b0;
    assign data[2624] = ~16'b0;
    assign data[2625] = ~16'b0;
    assign data[2626] = ~16'b0;
    assign data[2627] = ~16'b0;
    assign data[2628] = ~16'b0;
    assign data[2629] = ~16'b0;
    assign data[2630] = ~16'b0;
    assign data[2631] = ~16'b0;
    assign data[2632] = ~16'b0;
    assign data[2633] = ~16'b0;
    assign data[2634] = ~16'b0;
    assign data[2635] = ~16'b0;
    assign data[2636] = ~16'b0;
    assign data[2637] = ~16'b0;
    assign data[2638] = ~16'b0;
    assign data[2639] = ~16'b0;
    assign data[2640] = ~16'b0;
    assign data[2641] = ~16'b0;
    assign data[2642] = ~16'b0;
    assign data[2643] = ~16'b0;
    assign data[2644] = ~16'b0;
    assign data[2645] = ~16'b0;
    assign data[2646] = ~16'b0;
    assign data[2647] = ~16'b0;
    assign data[2648] = ~16'b0;
    assign data[2649] = ~16'b0;
    assign data[2650] = ~16'b0;
    assign data[2651] = ~16'b0;
    assign data[2652] = ~16'b0;
    assign data[2653] = ~16'b0;
    assign data[2654] = ~16'b0;
    assign data[2655] = ~16'b0;
    assign data[2656] = ~16'b0;
    assign data[2657] = ~16'b0;
    assign data[2658] = ~16'b0;
    assign data[2659] = ~16'b0;
    assign data[2660] = ~16'b0;
    assign data[2661] = ~16'b0;
    assign data[2662] = ~16'b0;
    assign data[2663] = ~16'b0;
    assign data[2664] = ~16'b0;
    assign data[2665] = ~16'b0;
    assign data[2666] = ~16'b0;
    assign data[2667] = ~16'b0;
    assign data[2668] = ~16'b0;
    assign data[2669] = ~16'b0;
    assign data[2670] = ~16'b0;
    assign data[2671] = ~16'b0;
    assign data[2672] = ~16'b0;
    assign data[2673] = ~16'b0;
    assign data[2674] = ~16'b0;
    assign data[2675] = ~16'b0;
    assign data[2676] = ~16'b0;
    assign data[2677] = ~16'b0;
    assign data[2678] = ~16'b0;
    assign data[2679] = ~16'b0;
    assign data[2680] = ~16'b0;
    assign data[2681] = ~16'b0;
    assign data[2682] = ~16'b0;
    assign data[2683] = ~16'b0;
    assign data[2684] = ~16'b0;
    assign data[2685] = ~16'b0;
    assign data[2686] = ~16'b0;
    assign data[2687] = ~16'b0;
    assign data[2688] = ~16'b0;
    assign data[2689] = ~16'b0;
    assign data[2690] = ~16'b0;
    assign data[2691] = ~16'b0;
    assign data[2692] = ~16'b0;
    assign data[2693] = ~16'b0;
    assign data[2694] = ~16'b0;
    assign data[2695] = ~16'b0;
    assign data[2696] = ~16'b0;
    assign data[2697] = ~16'b0;
    assign data[2698] = ~16'b0;
    assign data[2699] = ~16'b0;
    assign data[2700] = ~16'b0;
    assign data[2701] = ~16'b0;
    assign data[2702] = ~16'b0;
    assign data[2703] = ~16'b0;
    assign data[2704] = ~16'b0;
    assign data[2705] = ~16'b0;
    assign data[2706] = ~16'b0;
    assign data[2707] = ~16'b0;
    assign data[2708] = ~16'b0;
    assign data[2709] = ~16'b0;
    assign data[2710] = 16'b0;
    assign data[2711] = 16'b0;
    assign data[2712] = 16'b0;
    assign data[2713] = 16'b0;
    assign data[2714] = 16'b0;
    assign data[2715] = 16'b0;
    assign data[2716] = 16'b0;
    assign data[2717] = 16'b0;
    assign data[2718] = 16'b0;
    assign data[2719] = 16'b0;
    assign data[2720] = 16'b0;
    assign data[2721] = 16'b0;
    assign data[2722] = 16'b0;
    assign data[2723] = 16'b0;
    assign data[2724] = 16'b0;
    assign data[2725] = 16'b0;
    assign data[2726] = 16'b0;
    assign data[2727] = 16'b0;
    assign data[2728] = 16'b0;
    assign data[2729] = 16'b0;
    assign data[2730] = 16'b0;
    assign data[2731] = 16'b0;
    assign data[2732] = ~16'b0;
    assign data[2733] = ~16'b0;
    assign data[2734] = ~16'b0;
    assign data[2735] = ~16'b0;
    assign data[2736] = ~16'b0;
    assign data[2737] = ~16'b0;
    assign data[2738] = ~16'b0;
    assign data[2739] = ~16'b0;
    assign data[2740] = 16'b0;
    assign data[2741] = 16'b0;
    assign data[2742] = ~16'b0;
    assign data[2743] = ~16'b0;
    assign data[2744] = ~16'b0;
    assign data[2745] = ~16'b0;
    assign data[2746] = ~16'b0;
    assign data[2747] = ~16'b0;
    assign data[2748] = ~16'b0;
    assign data[2749] = ~16'b0;
    assign data[2750] = 16'b0;
    assign data[2751] = 16'b0;
    assign data[2752] = ~16'b0;
    assign data[2753] = ~16'b0;
    assign data[2754] = ~16'b0;
    assign data[2755] = ~16'b0;
    assign data[2756] = ~16'b0;
    assign data[2757] = ~16'b0;
    assign data[2758] = ~16'b0;
    assign data[2759] = ~16'b0;
    assign data[2760] = 16'b0;
    assign data[2761] = 16'b0;
    assign data[2762] = ~16'b0;
    assign data[2763] = ~16'b0;
    assign data[2764] = ~16'b0;
    assign data[2765] = ~16'b0;
    assign data[2766] = ~16'b0;
    assign data[2767] = ~16'b0;
    assign data[2768] = ~16'b0;
    assign data[2769] = ~16'b0;
    assign data[2770] = 16'b0;
    assign data[2771] = 16'b0;
    assign data[2772] = ~16'b0;
    assign data[2773] = ~16'b0;
    assign data[2774] = ~16'b0;
    assign data[2775] = ~16'b0;
    assign data[2776] = ~16'b0;
    assign data[2777] = ~16'b0;
    assign data[2778] = ~16'b0;
    assign data[2779] = ~16'b0;
    assign data[2780] = 16'b0;
    assign data[2781] = 16'b0;
    assign data[2782] = ~16'b0;
    assign data[2783] = ~16'b0;
    assign data[2784] = ~16'b0;
    assign data[2785] = ~16'b0;
    assign data[2786] = ~16'b0;
    assign data[2787] = ~16'b0;
    assign data[2788] = ~16'b0;
    assign data[2789] = ~16'b0;
    assign data[2790] = 16'b0;
    assign data[2791] = 16'b0;
    assign data[2792] = ~16'b0;
    assign data[2793] = ~16'b0;
    assign data[2794] = ~16'b0;
    assign data[2795] = ~16'b0;
    assign data[2796] = ~16'b0;
    assign data[2797] = ~16'b0;
    assign data[2798] = ~16'b0;
    assign data[2799] = ~16'b0;
    assign data[2800] = 16'b0;
    assign data[2801] = 16'b0;
    assign data[2802] = ~16'b0;
    assign data[2803] = ~16'b0;
    assign data[2804] = ~16'b0;
    assign data[2805] = ~16'b0;
    assign data[2806] = ~16'b0;
    assign data[2807] = ~16'b0;
    assign data[2808] = ~16'b0;
    assign data[2809] = ~16'b0;
    assign data[2810] = 16'b0;
    assign data[2811] = 16'b0;
    assign data[2812] = ~16'b0;
    assign data[2813] = ~16'b0;
    assign data[2814] = ~16'b0;
    assign data[2815] = ~16'b0;
    assign data[2816] = ~16'b0;
    assign data[2817] = ~16'b0;
    assign data[2818] = ~16'b0;
    assign data[2819] = ~16'b0;
    assign data[2820] = 16'b0;
    assign data[2821] = 16'b0;
    assign data[2822] = ~16'b0;
    assign data[2823] = ~16'b0;
    assign data[2824] = ~16'b0;
    assign data[2825] = ~16'b0;
    assign data[2826] = ~16'b0;
    assign data[2827] = ~16'b0;
    assign data[2828] = ~16'b0;
    assign data[2829] = ~16'b0;
    assign data[2830] = 16'b0;
    assign data[2831] = 16'b0;
    assign data[2832] = ~16'b0;
    assign data[2833] = ~16'b0;
    assign data[2834] = ~16'b0;
    assign data[2835] = ~16'b0;
    assign data[2836] = ~16'b0;
    assign data[2837] = ~16'b0;
    assign data[2838] = ~16'b0;
    assign data[2839] = ~16'b0;
    assign data[2840] = 16'b0;
    assign data[2841] = 16'b0;
    assign data[2842] = ~16'b0;
    assign data[2843] = ~16'b0;
    assign data[2844] = ~16'b0;
    assign data[2845] = ~16'b0;
    assign data[2846] = ~16'b0;
    assign data[2847] = ~16'b0;
    assign data[2848] = ~16'b0;
    assign data[2849] = ~16'b0;
    assign data[2850] = 16'b0;
    assign data[2851] = 16'b0;
    assign data[2852] = ~16'b0;
    assign data[2853] = ~16'b0;
    assign data[2854] = ~16'b0;
    assign data[2855] = ~16'b0;
    assign data[2856] = ~16'b0;
    assign data[2857] = ~16'b0;
    assign data[2858] = ~16'b0;
    assign data[2859] = ~16'b0;
    assign data[2860] = 16'b0;
    assign data[2861] = 16'b0;
    assign data[2862] = ~16'b0;
    assign data[2863] = ~16'b0;
    assign data[2864] = ~16'b0;
    assign data[2865] = ~16'b0;
    assign data[2866] = ~16'b0;
    assign data[2867] = ~16'b0;
    assign data[2868] = ~16'b0;
    assign data[2869] = ~16'b0;
    assign data[2870] = 16'b0;
    assign data[2871] = 16'b0;
    assign data[2872] = ~16'b0;
    assign data[2873] = ~16'b0;
    assign data[2874] = ~16'b0;
    assign data[2875] = ~16'b0;
    assign data[2876] = ~16'b0;
    assign data[2877] = ~16'b0;
    assign data[2878] = ~16'b0;
    assign data[2879] = ~16'b0;
    assign data[2880] = 16'b0;
    assign data[2881] = 16'b0;
    assign data[2882] = ~16'b0;
    assign data[2883] = ~16'b0;
    assign data[2884] = ~16'b0;
    assign data[2885] = ~16'b0;
    assign data[2886] = ~16'b0;
    assign data[2887] = ~16'b0;
    assign data[2888] = ~16'b0;
    assign data[2889] = ~16'b0;
    assign data[2890] = 16'b0;
    assign data[2891] = 16'b0;
    assign data[2892] = ~16'b0;
    assign data[2893] = ~16'b0;
    assign data[2894] = ~16'b0;
    assign data[2895] = ~16'b0;
    assign data[2896] = ~16'b0;
    assign data[2897] = ~16'b0;
    assign data[2898] = ~16'b0;
    assign data[2899] = ~16'b0;
    assign data[2900] = 16'b0;
    assign data[2901] = 16'b0;
    assign data[2902] = ~16'b0;
    assign data[2903] = ~16'b0;
    assign data[2904] = ~16'b0;
    assign data[2905] = ~16'b0;
    assign data[2906] = ~16'b0;
    assign data[2907] = ~16'b0;
    assign data[2908] = ~16'b0;
    assign data[2909] = ~16'b0;
    assign data[2910] = 16'b0;
    assign data[2911] = 16'b0;
    assign data[2912] = ~16'b0;
    assign data[2913] = ~16'b0;
    assign data[2914] = ~16'b0;
    assign data[2915] = ~16'b0;
    assign data[2916] = ~16'b0;
    assign data[2917] = ~16'b0;
    assign data[2918] = ~16'b0;
    assign data[2919] = ~16'b0;
    assign data[2920] = 16'b0;
    assign data[2921] = 16'b0;
    assign data[2922] = ~16'b0;
    assign data[2923] = ~16'b0;
    assign data[2924] = ~16'b0;
    assign data[2925] = ~16'b0;
    assign data[2926] = ~16'b0;
    assign data[2927] = ~16'b0;
    assign data[2928] = ~16'b0;
    assign data[2929] = ~16'b0;
    assign data[2930] = 16'b0;
    assign data[2931] = 16'b0;
    assign data[2932] = ~16'b0;
    assign data[2933] = ~16'b0;
    assign data[2934] = ~16'b0;
    assign data[2935] = ~16'b0;
    assign data[2936] = ~16'b0;
    assign data[2937] = ~16'b0;
    assign data[2938] = ~16'b0;
    assign data[2939] = ~16'b0;
    assign data[2940] = 16'b0;
    assign data[2941] = 16'b0;
    assign data[2942] = ~16'b0;
    assign data[2943] = ~16'b0;
    assign data[2944] = ~16'b0;
    assign data[2945] = ~16'b0;
    assign data[2946] = ~16'b0;
    assign data[2947] = ~16'b0;
    assign data[2948] = ~16'b0;
    assign data[2949] = ~16'b0;
    assign data[2950] = 16'b0;
    assign data[2951] = 16'b0;
    assign data[2952] = 16'b0;
    assign data[2953] = 16'b0;
    assign data[2954] = 16'b0;
    assign data[2955] = 16'b0;
    assign data[2956] = 16'b0;
    assign data[2957] = 16'b0;
    assign data[2958] = 16'b0;
    assign data[2959] = 16'b0;
    assign data[2960] = 16'b0;
    assign data[2961] = 16'b0;
    assign data[2962] = 16'b0;
    assign data[2963] = 16'b0;
    assign data[2964] = 16'b0;
    assign data[2965] = 16'b0;
    assign data[2966] = 16'b0;
    assign data[2967] = 16'b0;
    assign data[2968] = 16'b0;
    assign data[2969] = 16'b0;
    assign data[2970] = ~16'b0;
    assign data[2971] = ~16'b0;
    assign data[2972] = ~16'b0;
    assign data[2973] = ~16'b0;
    assign data[2974] = ~16'b0;
    assign data[2975] = ~16'b0;
    assign data[2976] = ~16'b0;
    assign data[2977] = ~16'b0;
    assign data[2978] = ~16'b0;
    assign data[2979] = ~16'b0;
    assign data[2980] = ~16'b0;
    assign data[2981] = ~16'b0;
    assign data[2982] = ~16'b0;
    assign data[2983] = ~16'b0;
    assign data[2984] = ~16'b0;
    assign data[2985] = ~16'b0;
    assign data[2986] = ~16'b0;
    assign data[2987] = ~16'b0;
    assign data[2988] = ~16'b0;
    assign data[2989] = ~16'b0;
    assign data[2990] = ~16'b0;
    assign data[2991] = ~16'b0;
    assign data[2992] = ~16'b0;
    assign data[2993] = ~16'b0;
    assign data[2994] = ~16'b0;
    assign data[2995] = ~16'b0;
    assign data[2996] = ~16'b0;
    assign data[2997] = ~16'b0;
    assign data[2998] = ~16'b0;
    assign data[2999] = ~16'b0;
    assign data[3000] = ~16'b0;
    assign data[3001] = ~16'b0;
    assign data[3002] = ~16'b0;
    assign data[3003] = ~16'b0;
    assign data[3004] = ~16'b0;
    assign data[3005] = ~16'b0;
    assign data[3006] = ~16'b0;
    assign data[3007] = ~16'b0;
    assign data[3008] = ~16'b0;
    assign data[3009] = ~16'b0;
    assign data[3010] = ~16'b0;
    assign data[3011] = ~16'b0;
    assign data[3012] = ~16'b0;
    assign data[3013] = ~16'b0;
    assign data[3014] = ~16'b0;
    assign data[3015] = ~16'b0;
    assign data[3016] = ~16'b0;
    assign data[3017] = ~16'b0;
    assign data[3018] = ~16'b0;
    assign data[3019] = ~16'b0;
    assign data[3020] = ~16'b0;
    assign data[3021] = ~16'b0;
    assign data[3022] = ~16'b0;
    assign data[3023] = ~16'b0;
    assign data[3024] = ~16'b0;
    assign data[3025] = ~16'b0;
    assign data[3026] = ~16'b0;
    assign data[3027] = ~16'b0;
    assign data[3028] = ~16'b0;
    assign data[3029] = ~16'b0;
    assign data[3030] = ~16'b0;
    assign data[3031] = ~16'b0;
    assign data[3032] = ~16'b0;
    assign data[3033] = ~16'b0;
    assign data[3034] = ~16'b0;
    assign data[3035] = ~16'b0;
    assign data[3036] = ~16'b0;
    assign data[3037] = ~16'b0;
    assign data[3038] = ~16'b0;
    assign data[3039] = ~16'b0;
    assign data[3040] = ~16'b0;
    assign data[3041] = ~16'b0;
    assign data[3042] = ~16'b0;
    assign data[3043] = ~16'b0;
    assign data[3044] = ~16'b0;
    assign data[3045] = ~16'b0;
    assign data[3046] = ~16'b0;
    assign data[3047] = ~16'b0;
    assign data[3048] = ~16'b0;
    assign data[3049] = ~16'b0;
    assign data[3050] = ~16'b0;
    assign data[3051] = ~16'b0;
    assign data[3052] = ~16'b0;
    assign data[3053] = ~16'b0;
    assign data[3054] = ~16'b0;
    assign data[3055] = ~16'b0;
    assign data[3056] = ~16'b0;
    assign data[3057] = ~16'b0;
    assign data[3058] = ~16'b0;
    assign data[3059] = ~16'b0;
    assign data[3060] = ~16'b0;
    assign data[3061] = ~16'b0;
    assign data[3062] = ~16'b0;
    assign data[3063] = ~16'b0;
    assign data[3064] = ~16'b0;
    assign data[3065] = ~16'b0;
    assign data[3066] = ~16'b0;
    assign data[3067] = ~16'b0;
    assign data[3068] = ~16'b0;
    assign data[3069] = ~16'b0;
    assign data[3070] = ~16'b0;
    assign data[3071] = ~16'b0;
    assign data[3072] = ~16'b0;
    assign data[3073] = ~16'b0;
    assign data[3074] = ~16'b0;
    assign data[3075] = ~16'b0;
    assign data[3076] = ~16'b0;
    assign data[3077] = ~16'b0;
    assign data[3078] = ~16'b0;
    assign data[3079] = ~16'b0;
    assign data[3080] = ~16'b0;
    assign data[3081] = ~16'b0;
    assign data[3082] = ~16'b0;
    assign data[3083] = ~16'b0;
    assign data[3084] = ~16'b0;
    assign data[3085] = ~16'b0;
    assign data[3086] = ~16'b0;
    assign data[3087] = ~16'b0;
    assign data[3088] = ~16'b0;
    assign data[3089] = ~16'b0;
    assign data[3090] = ~16'b0;
    assign data[3091] = ~16'b0;
    assign data[3092] = ~16'b0;
    assign data[3093] = ~16'b0;
    assign data[3094] = ~16'b0;
    assign data[3095] = ~16'b0;
    assign data[3096] = ~16'b0;
    assign data[3097] = ~16'b0;
    assign data[3098] = ~16'b0;
    assign data[3099] = ~16'b0;
    assign data[3100] = ~16'b0;
    assign data[3101] = ~16'b0;
    assign data[3102] = ~16'b0;
    assign data[3103] = ~16'b0;
    assign data[3104] = ~16'b0;
    assign data[3105] = ~16'b0;
    assign data[3106] = ~16'b0;
    assign data[3107] = ~16'b0;
    assign data[3108] = ~16'b0;
    assign data[3109] = ~16'b0;
    assign data[3110] = ~16'b0;
    assign data[3111] = ~16'b0;
    assign data[3112] = ~16'b0;
    assign data[3113] = ~16'b0;
    assign data[3114] = ~16'b0;
    assign data[3115] = ~16'b0;
    assign data[3116] = ~16'b0;
    assign data[3117] = ~16'b0;
    assign data[3118] = ~16'b0;
    assign data[3119] = ~16'b0;
    assign data[3120] = ~16'b0;
    assign data[3121] = ~16'b0;
    assign data[3122] = ~16'b0;
    assign data[3123] = ~16'b0;
    assign data[3124] = ~16'b0;
    assign data[3125] = ~16'b0;
    assign data[3126] = ~16'b0;
    assign data[3127] = ~16'b0;
    assign data[3128] = ~16'b0;
    assign data[3129] = ~16'b0;
    assign data[3130] = ~16'b0;
    assign data[3131] = ~16'b0;
    assign data[3132] = ~16'b0;
    assign data[3133] = ~16'b0;
    assign data[3134] = ~16'b0;
    assign data[3135] = ~16'b0;
    assign data[3136] = ~16'b0;
    assign data[3137] = ~16'b0;
    assign data[3138] = ~16'b0;
    assign data[3139] = ~16'b0;
    assign data[3140] = ~16'b0;
    assign data[3141] = ~16'b0;
    assign data[3142] = ~16'b0;
    assign data[3143] = ~16'b0;
    assign data[3144] = ~16'b0;
    assign data[3145] = ~16'b0;
    assign data[3146] = ~16'b0;
    assign data[3147] = ~16'b0;
    assign data[3148] = ~16'b0;
    assign data[3149] = ~16'b0;
    assign data[3150] = ~16'b0;
    assign data[3151] = ~16'b0;
    assign data[3152] = ~16'b0;
    assign data[3153] = ~16'b0;
    assign data[3154] = ~16'b0;
    assign data[3155] = ~16'b0;
    assign data[3156] = ~16'b0;
    assign data[3157] = ~16'b0;
    assign data[3158] = ~16'b0;
    assign data[3159] = ~16'b0;
    assign data[3160] = ~16'b0;
    assign data[3161] = ~16'b0;
    assign data[3162] = ~16'b0;
    assign data[3163] = ~16'b0;
    assign data[3164] = ~16'b0;
    assign data[3165] = ~16'b0;
    assign data[3166] = ~16'b0;
    assign data[3167] = ~16'b0;
    assign data[3168] = ~16'b0;
    assign data[3169] = ~16'b0;
    assign data[3170] = ~16'b0;
    assign data[3171] = ~16'b0;
    assign data[3172] = ~16'b0;
    assign data[3173] = ~16'b0;
    assign data[3174] = ~16'b0;
    assign data[3175] = ~16'b0;
    assign data[3176] = ~16'b0;
    assign data[3177] = ~16'b0;
    assign data[3178] = ~16'b0;
    assign data[3179] = ~16'b0;
    assign data[3180] = ~16'b0;
    assign data[3181] = ~16'b0;
    assign data[3182] = ~16'b0;
    assign data[3183] = ~16'b0;
    assign data[3184] = ~16'b0;
    assign data[3185] = ~16'b0;
    assign data[3186] = ~16'b0;
    assign data[3187] = ~16'b0;
    assign data[3188] = ~16'b0;
    assign data[3189] = ~16'b0;
    assign data[3190] = ~16'b0;
    assign data[3191] = ~16'b0;
    assign data[3192] = ~16'b0;
    assign data[3193] = ~16'b0;
    assign data[3194] = ~16'b0;
    assign data[3195] = ~16'b0;
    assign data[3196] = ~16'b0;
    assign data[3197] = ~16'b0;
    assign data[3198] = ~16'b0;
    assign data[3199] = ~16'b0;
    assign data[3200] = ~16'b0;
    assign data[3201] = ~16'b0;
    assign data[3202] = ~16'b0;
    assign data[3203] = ~16'b0;
    assign data[3204] = ~16'b0;
    assign data[3205] = ~16'b0;
    assign data[3206] = ~16'b0;
    assign data[3207] = ~16'b0;
    assign data[3208] = ~16'b0;
    assign data[3209] = ~16'b0;
    assign data[3210] = ~16'b0;
    assign data[3211] = ~16'b0;
    assign data[3212] = ~16'b0;
    assign data[3213] = ~16'b0;
    assign data[3214] = ~16'b0;
    assign data[3215] = ~16'b0;
    assign data[3216] = ~16'b0;
    assign data[3217] = ~16'b0;
    assign data[3218] = ~16'b0;
    assign data[3219] = ~16'b0;
    assign data[3220] = ~16'b0;
    assign data[3221] = ~16'b0;
    assign data[3222] = ~16'b0;
    assign data[3223] = ~16'b0;
    assign data[3224] = ~16'b0;
    assign data[3225] = ~16'b0;
    assign data[3226] = ~16'b0;
    assign data[3227] = ~16'b0;
    assign data[3228] = ~16'b0;
    assign data[3229] = ~16'b0;
    assign data[3230] = ~16'b0;
    assign data[3231] = ~16'b0;
    assign data[3232] = ~16'b0;
    assign data[3233] = ~16'b0;
    assign data[3234] = ~16'b0;
    assign data[3235] = ~16'b0;
    assign data[3236] = ~16'b0;
    assign data[3237] = ~16'b0;
    assign data[3238] = ~16'b0;
    assign data[3239] = ~16'b0;
    assign data[3240] = ~16'b0;
    assign data[3241] = ~16'b0;
    assign data[3242] = ~16'b0;
    assign data[3243] = ~16'b0;
    assign data[3244] = ~16'b0;
    assign data[3245] = ~16'b0;
    assign data[3246] = ~16'b0;
    assign data[3247] = ~16'b0;
    assign data[3248] = ~16'b0;
    assign data[3249] = ~16'b0;
    assign data[3250] = ~16'b0;
    assign data[3251] = ~16'b0;
    assign data[3252] = ~16'b0;
    assign data[3253] = ~16'b0;
    assign data[3254] = ~16'b0;
    assign data[3255] = ~16'b0;
    assign data[3256] = ~16'b0;
    assign data[3257] = ~16'b0;
    assign data[3258] = ~16'b0;
    assign data[3259] = ~16'b0;
    assign data[3260] = ~16'b0;
    assign data[3261] = ~16'b0;
    assign data[3262] = ~16'b0;
    assign data[3263] = ~16'b0;
    assign data[3264] = ~16'b0;
    assign data[3265] = ~16'b0;
    assign data[3266] = ~16'b0;
    assign data[3267] = ~16'b0;
    assign data[3268] = ~16'b0;
    assign data[3269] = ~16'b0;
    assign data[3270] = ~16'b0;
    assign data[3271] = ~16'b0;
    assign data[3272] = ~16'b0;
    assign data[3273] = ~16'b0;
    assign data[3274] = ~16'b0;
    assign data[3275] = ~16'b0;
    assign data[3276] = ~16'b0;
    assign data[3277] = ~16'b0;
    assign data[3278] = ~16'b0;
    assign data[3279] = ~16'b0;
    assign data[3280] = ~16'b0;
    assign data[3281] = ~16'b0;
    assign data[3282] = ~16'b0;
    assign data[3283] = ~16'b0;
    assign data[3284] = ~16'b0;
    assign data[3285] = ~16'b0;
    assign data[3286] = ~16'b0;
    assign data[3287] = ~16'b0;
    assign data[3288] = ~16'b0;
    assign data[3289] = ~16'b0;
    assign data[3290] = 16'b0;
    assign data[3291] = 16'b0;
    assign data[3292] = 16'b0;
    assign data[3293] = 16'b0;
    assign data[3294] = 16'b0;
    assign data[3295] = 16'b0;
    assign data[3296] = 16'b0;
    assign data[3297] = 16'b0;
    assign data[3298] = 16'b0;
    assign data[3299] = 16'b0;
    assign data[3300] = 16'b0;
    assign data[3301] = 16'b0;
    assign data[3302] = 16'b0;
    assign data[3303] = 16'b0;
    assign data[3304] = 16'b0;
    assign data[3305] = 16'b0;
    assign data[3306] = 16'b0;
    assign data[3307] = 16'b0;
    assign data[3308] = 16'b0;
    assign data[3309] = 16'b0;
    assign data[3310] = 16'b0;
    assign data[3311] = 16'b0;
    assign data[3312] = ~16'b0;
    assign data[3313] = ~16'b0;
    assign data[3314] = ~16'b0;
    assign data[3315] = ~16'b0;
    assign data[3316] = ~16'b0;
    assign data[3317] = ~16'b0;
    assign data[3318] = ~16'b0;
    assign data[3319] = ~16'b0;
    assign data[3320] = 16'b0;
    assign data[3321] = 16'b0;
    assign data[3322] = ~16'b0;
    assign data[3323] = ~16'b0;
    assign data[3324] = ~16'b0;
    assign data[3325] = ~16'b0;
    assign data[3326] = ~16'b0;
    assign data[3327] = ~16'b0;
    assign data[3328] = ~16'b0;
    assign data[3329] = ~16'b0;
    assign data[3330] = 16'b0;
    assign data[3331] = 16'b0;
    assign data[3332] = ~16'b0;
    assign data[3333] = ~16'b0;
    assign data[3334] = ~16'b0;
    assign data[3335] = ~16'b0;
    assign data[3336] = ~16'b0;
    assign data[3337] = ~16'b0;
    assign data[3338] = ~16'b0;
    assign data[3339] = ~16'b0;
    assign data[3340] = 16'b0;
    assign data[3341] = 16'b0;
    assign data[3342] = ~16'b0;
    assign data[3343] = ~16'b0;
    assign data[3344] = ~16'b0;
    assign data[3345] = ~16'b0;
    assign data[3346] = ~16'b0;
    assign data[3347] = ~16'b0;
    assign data[3348] = ~16'b0;
    assign data[3349] = ~16'b0;
    assign data[3350] = 16'b0;
    assign data[3351] = 16'b0;
    assign data[3352] = ~16'b0;
    assign data[3353] = ~16'b0;
    assign data[3354] = ~16'b0;
    assign data[3355] = ~16'b0;
    assign data[3356] = ~16'b0;
    assign data[3357] = ~16'b0;
    assign data[3358] = ~16'b0;
    assign data[3359] = ~16'b0;
    assign data[3360] = 16'b0;
    assign data[3361] = 16'b0;
    assign data[3362] = ~16'b0;
    assign data[3363] = ~16'b0;
    assign data[3364] = ~16'b0;
    assign data[3365] = ~16'b0;
    assign data[3366] = ~16'b0;
    assign data[3367] = ~16'b0;
    assign data[3368] = ~16'b0;
    assign data[3369] = ~16'b0;
    assign data[3370] = 16'b0;
    assign data[3371] = 16'b0;
    assign data[3372] = ~16'b0;
    assign data[3373] = ~16'b0;
    assign data[3374] = ~16'b0;
    assign data[3375] = ~16'b0;
    assign data[3376] = ~16'b0;
    assign data[3377] = ~16'b0;
    assign data[3378] = ~16'b0;
    assign data[3379] = ~16'b0;
    assign data[3380] = 16'b0;
    assign data[3381] = 16'b0;
    assign data[3382] = ~16'b0;
    assign data[3383] = ~16'b0;
    assign data[3384] = ~16'b0;
    assign data[3385] = ~16'b0;
    assign data[3386] = ~16'b0;
    assign data[3387] = ~16'b0;
    assign data[3388] = ~16'b0;
    assign data[3389] = ~16'b0;
    assign data[3390] = 16'b0;
    assign data[3391] = 16'b0;
    assign data[3392] = ~16'b0;
    assign data[3393] = ~16'b0;
    assign data[3394] = ~16'b0;
    assign data[3395] = ~16'b0;
    assign data[3396] = ~16'b0;
    assign data[3397] = ~16'b0;
    assign data[3398] = ~16'b0;
    assign data[3399] = ~16'b0;
    assign data[3400] = 16'b0;
    assign data[3401] = 16'b0;
    assign data[3402] = ~16'b0;
    assign data[3403] = ~16'b0;
    assign data[3404] = ~16'b0;
    assign data[3405] = ~16'b0;
    assign data[3406] = ~16'b0;
    assign data[3407] = ~16'b0;
    assign data[3408] = ~16'b0;
    assign data[3409] = ~16'b0;
    assign data[3410] = 16'b0;
    assign data[3411] = 16'b0;
    assign data[3412] = ~16'b0;
    assign data[3413] = ~16'b0;
    assign data[3414] = ~16'b0;
    assign data[3415] = ~16'b0;
    assign data[3416] = ~16'b0;
    assign data[3417] = ~16'b0;
    assign data[3418] = ~16'b0;
    assign data[3419] = ~16'b0;
    assign data[3420] = 16'b0;
    assign data[3421] = 16'b0;
    assign data[3422] = ~16'b0;
    assign data[3423] = ~16'b0;
    assign data[3424] = ~16'b0;
    assign data[3425] = ~16'b0;
    assign data[3426] = ~16'b0;
    assign data[3427] = ~16'b0;
    assign data[3428] = ~16'b0;
    assign data[3429] = ~16'b0;
    assign data[3430] = 16'b0;
    assign data[3431] = 16'b0;
    assign data[3432] = ~16'b0;
    assign data[3433] = ~16'b0;
    assign data[3434] = ~16'b0;
    assign data[3435] = ~16'b0;
    assign data[3436] = ~16'b0;
    assign data[3437] = ~16'b0;
    assign data[3438] = ~16'b0;
    assign data[3439] = ~16'b0;
    assign data[3440] = 16'b0;
    assign data[3441] = 16'b0;
    assign data[3442] = ~16'b0;
    assign data[3443] = ~16'b0;
    assign data[3444] = ~16'b0;
    assign data[3445] = ~16'b0;
    assign data[3446] = ~16'b0;
    assign data[3447] = ~16'b0;
    assign data[3448] = ~16'b0;
    assign data[3449] = ~16'b0;
    assign data[3450] = 16'b0;
    assign data[3451] = 16'b0;
    assign data[3452] = ~16'b0;
    assign data[3453] = ~16'b0;
    assign data[3454] = ~16'b0;
    assign data[3455] = ~16'b0;
    assign data[3456] = ~16'b0;
    assign data[3457] = ~16'b0;
    assign data[3458] = ~16'b0;
    assign data[3459] = ~16'b0;
    assign data[3460] = 16'b0;
    assign data[3461] = 16'b0;
    assign data[3462] = ~16'b0;
    assign data[3463] = ~16'b0;
    assign data[3464] = ~16'b0;
    assign data[3465] = ~16'b0;
    assign data[3466] = ~16'b0;
    assign data[3467] = ~16'b0;
    assign data[3468] = ~16'b0;
    assign data[3469] = ~16'b0;
    assign data[3470] = 16'b0;
    assign data[3471] = 16'b0;
    assign data[3472] = ~16'b0;
    assign data[3473] = ~16'b0;
    assign data[3474] = ~16'b0;
    assign data[3475] = ~16'b0;
    assign data[3476] = ~16'b0;
    assign data[3477] = ~16'b0;
    assign data[3478] = ~16'b0;
    assign data[3479] = ~16'b0;
    assign data[3480] = 16'b0;
    assign data[3481] = 16'b0;
    assign data[3482] = ~16'b0;
    assign data[3483] = ~16'b0;
    assign data[3484] = ~16'b0;
    assign data[3485] = ~16'b0;
    assign data[3486] = ~16'b0;
    assign data[3487] = ~16'b0;
    assign data[3488] = ~16'b0;
    assign data[3489] = ~16'b0;
    assign data[3490] = 16'b0;
    assign data[3491] = 16'b0;
    assign data[3492] = ~16'b0;
    assign data[3493] = ~16'b0;
    assign data[3494] = ~16'b0;
    assign data[3495] = ~16'b0;
    assign data[3496] = ~16'b0;
    assign data[3497] = ~16'b0;
    assign data[3498] = ~16'b0;
    assign data[3499] = ~16'b0;
    assign data[3500] = 16'b0;
    assign data[3501] = 16'b0;
    assign data[3502] = ~16'b0;
    assign data[3503] = ~16'b0;
    assign data[3504] = ~16'b0;
    assign data[3505] = ~16'b0;
    assign data[3506] = ~16'b0;
    assign data[3507] = ~16'b0;
    assign data[3508] = ~16'b0;
    assign data[3509] = ~16'b0;
    assign data[3510] = 16'b0;
    assign data[3511] = 16'b0;
    assign data[3512] = ~16'b0;
    assign data[3513] = ~16'b0;
    assign data[3514] = ~16'b0;
    assign data[3515] = ~16'b0;
    assign data[3516] = ~16'b0;
    assign data[3517] = ~16'b0;
    assign data[3518] = ~16'b0;
    assign data[3519] = ~16'b0;
    assign data[3520] = 16'b0;
    assign data[3521] = 16'b0;
    assign data[3522] = ~16'b0;
    assign data[3523] = ~16'b0;
    assign data[3524] = ~16'b0;
    assign data[3525] = ~16'b0;
    assign data[3526] = ~16'b0;
    assign data[3527] = ~16'b0;
    assign data[3528] = ~16'b0;
    assign data[3529] = ~16'b0;
    assign data[3530] = 16'b0;
    assign data[3531] = 16'b0;
    assign data[3532] = ~16'b0;
    assign data[3533] = ~16'b0;
    assign data[3534] = ~16'b0;
    assign data[3535] = ~16'b0;
    assign data[3536] = ~16'b0;
    assign data[3537] = ~16'b0;
    assign data[3538] = ~16'b0;
    assign data[3539] = ~16'b0;
    assign data[3540] = 16'b0;
    assign data[3541] = 16'b0;
    assign data[3542] = ~16'b0;
    assign data[3543] = ~16'b0;
    assign data[3544] = ~16'b0;
    assign data[3545] = ~16'b0;
    assign data[3546] = ~16'b0;
    assign data[3547] = ~16'b0;
    assign data[3548] = ~16'b0;
    assign data[3549] = ~16'b0;
    assign data[3550] = 16'b0;
    assign data[3551] = 16'b0;
    assign data[3552] = ~16'b0;
    assign data[3553] = ~16'b0;
    assign data[3554] = ~16'b0;
    assign data[3555] = ~16'b0;
    assign data[3556] = ~16'b0;
    assign data[3557] = ~16'b0;
    assign data[3558] = ~16'b0;
    assign data[3559] = ~16'b0;
    assign data[3560] = 16'b0;
    assign data[3561] = 16'b0;
    assign data[3562] = ~16'b0;
    assign data[3563] = ~16'b0;
    assign data[3564] = ~16'b0;
    assign data[3565] = ~16'b0;
    assign data[3566] = ~16'b0;
    assign data[3567] = ~16'b0;
    assign data[3568] = ~16'b0;
    assign data[3569] = ~16'b0;
    assign data[3570] = 16'b0;
    assign data[3571] = 16'b0;
    assign data[3572] = ~16'b0;
    assign data[3573] = ~16'b0;
    assign data[3574] = ~16'b0;
    assign data[3575] = ~16'b0;
    assign data[3576] = ~16'b0;
    assign data[3577] = ~16'b0;
    assign data[3578] = ~16'b0;
    assign data[3579] = ~16'b0;
    assign data[3580] = 16'b0;
    assign data[3581] = 16'b0;
    assign data[3582] = ~16'b0;
    assign data[3583] = ~16'b0;
    assign data[3584] = ~16'b0;
    assign data[3585] = ~16'b0;
    assign data[3586] = ~16'b0;
    assign data[3587] = ~16'b0;
    assign data[3588] = ~16'b0;
    assign data[3589] = ~16'b0;
    assign data[3590] = 16'b0;
    assign data[3591] = 16'b0;
    assign data[3592] = ~16'b0;
    assign data[3593] = ~16'b0;
    assign data[3594] = ~16'b0;
    assign data[3595] = ~16'b0;
    assign data[3596] = ~16'b0;
    assign data[3597] = ~16'b0;
    assign data[3598] = ~16'b0;
    assign data[3599] = ~16'b0;
    assign data[3600] = 16'b0;
    assign data[3601] = 16'b0;
    assign data[3602] = ~16'b0;
    assign data[3603] = ~16'b0;
    assign data[3604] = ~16'b0;
    assign data[3605] = ~16'b0;
    assign data[3606] = ~16'b0;
    assign data[3607] = ~16'b0;
    assign data[3608] = ~16'b0;
    assign data[3609] = ~16'b0;
    assign data[3610] = 16'b0;
    assign data[3611] = 16'b0;
    assign data[3612] = ~16'b0;
    assign data[3613] = ~16'b0;
    assign data[3614] = ~16'b0;
    assign data[3615] = ~16'b0;
    assign data[3616] = ~16'b0;
    assign data[3617] = ~16'b0;
    assign data[3618] = ~16'b0;
    assign data[3619] = ~16'b0;
    assign data[3620] = 16'b0;
    assign data[3621] = 16'b0;
    assign data[3622] = ~16'b0;
    assign data[3623] = ~16'b0;
    assign data[3624] = ~16'b0;
    assign data[3625] = ~16'b0;
    assign data[3626] = ~16'b0;
    assign data[3627] = ~16'b0;
    assign data[3628] = ~16'b0;
    assign data[3629] = ~16'b0;
    assign data[3630] = 16'b0;
    assign data[3631] = 16'b0;
    assign data[3632] = ~16'b0;
    assign data[3633] = ~16'b0;
    assign data[3634] = ~16'b0;
    assign data[3635] = ~16'b0;
    assign data[3636] = ~16'b0;
    assign data[3637] = ~16'b0;
    assign data[3638] = ~16'b0;
    assign data[3639] = ~16'b0;
    assign data[3640] = 16'b0;
    assign data[3641] = 16'b0;
    assign data[3642] = ~16'b0;
    assign data[3643] = ~16'b0;
    assign data[3644] = ~16'b0;
    assign data[3645] = ~16'b0;
    assign data[3646] = ~16'b0;
    assign data[3647] = ~16'b0;
    assign data[3648] = ~16'b0;
    assign data[3649] = ~16'b0;
    assign data[3650] = 16'b0;
    assign data[3651] = 16'b0;
    assign data[3652] = ~16'b0;
    assign data[3653] = ~16'b0;
    assign data[3654] = ~16'b0;
    assign data[3655] = ~16'b0;
    assign data[3656] = ~16'b0;
    assign data[3657] = ~16'b0;
    assign data[3658] = ~16'b0;
    assign data[3659] = ~16'b0;
    assign data[3660] = 16'b0;
    assign data[3661] = 16'b0;
    assign data[3662] = ~16'b0;
    assign data[3663] = ~16'b0;
    assign data[3664] = ~16'b0;
    assign data[3665] = ~16'b0;
    assign data[3666] = ~16'b0;
    assign data[3667] = ~16'b0;
    assign data[3668] = ~16'b0;
    assign data[3669] = ~16'b0;
    assign data[3670] = 16'b0;
    assign data[3671] = 16'b0;
    assign data[3672] = ~16'b0;
    assign data[3673] = ~16'b0;
    assign data[3674] = ~16'b0;
    assign data[3675] = ~16'b0;
    assign data[3676] = ~16'b0;
    assign data[3677] = ~16'b0;
    assign data[3678] = ~16'b0;
    assign data[3679] = ~16'b0;
    assign data[3680] = 16'b0;
    assign data[3681] = 16'b0;
    assign data[3682] = ~16'b0;
    assign data[3683] = ~16'b0;
    assign data[3684] = ~16'b0;
    assign data[3685] = ~16'b0;
    assign data[3686] = ~16'b0;
    assign data[3687] = ~16'b0;
    assign data[3688] = ~16'b0;
    assign data[3689] = ~16'b0;
    assign data[3690] = 16'b0;
    assign data[3691] = 16'b0;
    assign data[3692] = ~16'b0;
    assign data[3693] = ~16'b0;
    assign data[3694] = ~16'b0;
    assign data[3695] = ~16'b0;
    assign data[3696] = ~16'b0;
    assign data[3697] = ~16'b0;
    assign data[3698] = ~16'b0;
    assign data[3699] = ~16'b0;
    assign data[3700] = 16'b0;
    assign data[3701] = 16'b0;
    assign data[3702] = ~16'b0;
    assign data[3703] = ~16'b0;
    assign data[3704] = ~16'b0;
    assign data[3705] = ~16'b0;
    assign data[3706] = ~16'b0;
    assign data[3707] = ~16'b0;
    assign data[3708] = ~16'b0;
    assign data[3709] = ~16'b0;
    assign data[3710] = 16'b0;
    assign data[3711] = 16'b0;
    assign data[3712] = ~16'b0;
    assign data[3713] = ~16'b0;
    assign data[3714] = ~16'b0;
    assign data[3715] = ~16'b0;
    assign data[3716] = ~16'b0;
    assign data[3717] = ~16'b0;
    assign data[3718] = ~16'b0;
    assign data[3719] = ~16'b0;
    assign data[3720] = 16'b0;
    assign data[3721] = 16'b0;
    assign data[3722] = ~16'b0;
    assign data[3723] = ~16'b0;
    assign data[3724] = ~16'b0;
    assign data[3725] = ~16'b0;
    assign data[3726] = ~16'b0;
    assign data[3727] = ~16'b0;
    assign data[3728] = ~16'b0;
    assign data[3729] = ~16'b0;
    assign data[3730] = 16'b0;
    assign data[3731] = 16'b0;
    assign data[3732] = ~16'b0;
    assign data[3733] = ~16'b0;
    assign data[3734] = ~16'b0;
    assign data[3735] = ~16'b0;
    assign data[3736] = ~16'b0;
    assign data[3737] = ~16'b0;
    assign data[3738] = ~16'b0;
    assign data[3739] = ~16'b0;
    assign data[3740] = 16'b0;
    assign data[3741] = 16'b0;
    assign data[3742] = ~16'b0;
    assign data[3743] = ~16'b0;
    assign data[3744] = ~16'b0;
    assign data[3745] = ~16'b0;
    assign data[3746] = ~16'b0;
    assign data[3747] = ~16'b0;
    assign data[3748] = ~16'b0;
    assign data[3749] = ~16'b0;
    assign data[3750] = 16'b0;
    assign data[3751] = 16'b0;
    assign data[3752] = ~16'b0;
    assign data[3753] = ~16'b0;
    assign data[3754] = ~16'b0;
    assign data[3755] = ~16'b0;
    assign data[3756] = ~16'b0;
    assign data[3757] = ~16'b0;
    assign data[3758] = ~16'b0;
    assign data[3759] = ~16'b0;
    assign data[3760] = 16'b0;
    assign data[3761] = 16'b0;
    assign data[3762] = ~16'b0;
    assign data[3763] = ~16'b0;
    assign data[3764] = ~16'b0;
    assign data[3765] = ~16'b0;
    assign data[3766] = ~16'b0;
    assign data[3767] = ~16'b0;
    assign data[3768] = ~16'b0;
    assign data[3769] = ~16'b0;
    assign data[3770] = 16'b0;
    assign data[3771] = 16'b0;
    assign data[3772] = 16'b0;
    assign data[3773] = 16'b0;
    assign data[3774] = 16'b0;
    assign data[3775] = 16'b0;
    assign data[3776] = 16'b0;
    assign data[3777] = 16'b0;
    assign data[3778] = 16'b0;
    assign data[3779] = 16'b0;
    assign data[3780] = 16'b0;
    assign data[3781] = 16'b0;
    assign data[3782] = 16'b0;
    assign data[3783] = 16'b0;
    assign data[3784] = 16'b0;
    assign data[3785] = 16'b0;
    assign data[3786] = 16'b0;
    assign data[3787] = 16'b0;
    assign data[3788] = 16'b0;
    assign data[3789] = 16'b0;
    assign data[3790] = ~16'b0;
    assign data[3791] = ~16'b0;
    assign data[3792] = ~16'b0;
    assign data[3793] = ~16'b0;
    assign data[3794] = ~16'b0;
    assign data[3795] = ~16'b0;
    assign data[3796] = ~16'b0;
    assign data[3797] = ~16'b0;
    assign data[3798] = ~16'b0;
    assign data[3799] = ~16'b0;
    assign data[3800] = ~16'b0;
    assign data[3801] = ~16'b0;
    assign data[3802] = ~16'b0;
    assign data[3803] = ~16'b0;
    assign data[3804] = ~16'b0;
    assign data[3805] = ~16'b0;
    assign data[3806] = ~16'b0;
    assign data[3807] = ~16'b0;
    assign data[3808] = ~16'b0;
    assign data[3809] = ~16'b0;
    assign data[3810] = ~16'b0;
    assign data[3811] = ~16'b0;
    assign data[3812] = ~16'b0;
    assign data[3813] = ~16'b0;
    assign data[3814] = ~16'b0;
    assign data[3815] = ~16'b0;
    assign data[3816] = ~16'b0;
    assign data[3817] = ~16'b0;
    assign data[3818] = ~16'b0;
    assign data[3819] = ~16'b0;
    assign data[3820] = ~16'b0;
    assign data[3821] = ~16'b0;
    assign data[3822] = ~16'b0;
    assign data[3823] = ~16'b0;
    assign data[3824] = ~16'b0;
    assign data[3825] = ~16'b0;
    assign data[3826] = ~16'b0;
    assign data[3827] = ~16'b0;
    assign data[3828] = ~16'b0;
    assign data[3829] = ~16'b0;
    assign data[3830] = ~16'b0;
    assign data[3831] = ~16'b0;
    assign data[3832] = ~16'b0;
    assign data[3833] = ~16'b0;
    assign data[3834] = ~16'b0;
    assign data[3835] = ~16'b0;
    assign data[3836] = ~16'b0;
    assign data[3837] = ~16'b0;
    assign data[3838] = ~16'b0;
    assign data[3839] = ~16'b0;
    assign data[3840] = ~16'b0;
    assign data[3841] = ~16'b0;
    assign data[3842] = ~16'b0;
    assign data[3843] = ~16'b0;
    assign data[3844] = ~16'b0;
    assign data[3845] = ~16'b0;
    assign data[3846] = ~16'b0;
    assign data[3847] = ~16'b0;
    assign data[3848] = ~16'b0;
    assign data[3849] = ~16'b0;
    assign data[3850] = ~16'b0;
    assign data[3851] = ~16'b0;
    assign data[3852] = ~16'b0;
    assign data[3853] = ~16'b0;
    assign data[3854] = ~16'b0;
    assign data[3855] = ~16'b0;
    assign data[3856] = ~16'b0;
    assign data[3857] = ~16'b0;
    assign data[3858] = ~16'b0;
    assign data[3859] = ~16'b0;
    assign data[3860] = ~16'b0;
    assign data[3861] = ~16'b0;
    assign data[3862] = ~16'b0;
    assign data[3863] = ~16'b0;
    assign data[3864] = ~16'b0;
    assign data[3865] = ~16'b0;
    assign data[3866] = ~16'b0;
    assign data[3867] = ~16'b0;
    assign data[3868] = ~16'b0;
    assign data[3869] = ~16'b0;
    assign data[3870] = ~16'b0;
    assign data[3871] = ~16'b0;
    assign data[3872] = ~16'b0;
    assign data[3873] = ~16'b0;
    assign data[3874] = ~16'b0;
    assign data[3875] = ~16'b0;
    assign data[3876] = ~16'b0;
    assign data[3877] = ~16'b0;
    assign data[3878] = ~16'b0;
    assign data[3879] = ~16'b0;
    assign data[3880] = ~16'b0;
    assign data[3881] = ~16'b0;
    assign data[3882] = ~16'b0;
    assign data[3883] = ~16'b0;
    assign data[3884] = ~16'b0;
    assign data[3885] = ~16'b0;
    assign data[3886] = ~16'b0;
    assign data[3887] = ~16'b0;
    assign data[3888] = ~16'b0;
    assign data[3889] = ~16'b0;
    assign data[3890] = ~16'b0;
    assign data[3891] = ~16'b0;
    assign data[3892] = ~16'b0;
    assign data[3893] = ~16'b0;
    assign data[3894] = ~16'b0;
    assign data[3895] = ~16'b0;
    assign data[3896] = ~16'b0;
    assign data[3897] = ~16'b0;
    assign data[3898] = ~16'b0;
    assign data[3899] = ~16'b0;
    assign data[3900] = ~16'b0;
    assign data[3901] = ~16'b0;
    assign data[3902] = ~16'b0;
    assign data[3903] = ~16'b0;
    assign data[3904] = ~16'b0;
    assign data[3905] = ~16'b0;
    assign data[3906] = ~16'b0;
    assign data[3907] = ~16'b0;
    assign data[3908] = ~16'b0;
    assign data[3909] = ~16'b0;
    assign data[3910] = ~16'b0;
    assign data[3911] = ~16'b0;
    assign data[3912] = ~16'b0;
    assign data[3913] = ~16'b0;
    assign data[3914] = ~16'b0;
    assign data[3915] = ~16'b0;
    assign data[3916] = ~16'b0;
    assign data[3917] = ~16'b0;
    assign data[3918] = ~16'b0;
    assign data[3919] = ~16'b0;
    assign data[3920] = ~16'b0;
    assign data[3921] = ~16'b0;
    assign data[3922] = ~16'b0;
    assign data[3923] = ~16'b0;
    assign data[3924] = ~16'b0;
    assign data[3925] = ~16'b0;
    assign data[3926] = ~16'b0;
    assign data[3927] = ~16'b0;
    assign data[3928] = ~16'b0;
    assign data[3929] = ~16'b0;
    assign data[3930] = ~16'b0;
    assign data[3931] = ~16'b0;
    assign data[3932] = ~16'b0;
    assign data[3933] = ~16'b0;
    assign data[3934] = ~16'b0;
    assign data[3935] = ~16'b0;
    assign data[3936] = ~16'b0;
    assign data[3937] = ~16'b0;
    assign data[3938] = ~16'b0;
    assign data[3939] = ~16'b0;
    assign data[3940] = ~16'b0;
    assign data[3941] = ~16'b0;
    assign data[3942] = ~16'b0;
    assign data[3943] = ~16'b0;
    assign data[3944] = ~16'b0;
    assign data[3945] = ~16'b0;
    assign data[3946] = ~16'b0;
    assign data[3947] = ~16'b0;
    assign data[3948] = ~16'b0;
    assign data[3949] = ~16'b0;
    assign data[3950] = ~16'b0;
    assign data[3951] = ~16'b0;
    assign data[3952] = ~16'b0;
    assign data[3953] = ~16'b0;
    assign data[3954] = ~16'b0;
    assign data[3955] = ~16'b0;
    assign data[3956] = ~16'b0;
    assign data[3957] = ~16'b0;
    assign data[3958] = ~16'b0;
    assign data[3959] = ~16'b0;
    assign data[3960] = ~16'b0;
    assign data[3961] = ~16'b0;
    assign data[3962] = ~16'b0;
    assign data[3963] = ~16'b0;
    assign data[3964] = ~16'b0;
    assign data[3965] = ~16'b0;
    assign data[3966] = ~16'b0;
    assign data[3967] = ~16'b0;
    assign data[3968] = ~16'b0;
    assign data[3969] = ~16'b0;
    assign data[3970] = ~16'b0;
    assign data[3971] = ~16'b0;
    assign data[3972] = ~16'b0;
    assign data[3973] = ~16'b0;
    assign data[3974] = ~16'b0;
    assign data[3975] = ~16'b0;
    assign data[3976] = ~16'b0;
    assign data[3977] = ~16'b0;
    assign data[3978] = ~16'b0;
    assign data[3979] = ~16'b0;
    assign data[3980] = ~16'b0;
    assign data[3981] = ~16'b0;
    assign data[3982] = ~16'b0;
    assign data[3983] = ~16'b0;
    assign data[3984] = ~16'b0;
    assign data[3985] = ~16'b0;
    assign data[3986] = ~16'b0;
    assign data[3987] = ~16'b0;
    assign data[3988] = ~16'b0;
    assign data[3989] = ~16'b0;
    assign data[3990] = ~16'b0;
    assign data[3991] = ~16'b0;
    assign data[3992] = ~16'b0;
    assign data[3993] = ~16'b0;
    assign data[3994] = ~16'b0;
    assign data[3995] = ~16'b0;
    assign data[3996] = ~16'b0;
    assign data[3997] = ~16'b0;
    assign data[3998] = ~16'b0;
    assign data[3999] = ~16'b0;
    assign data[4000] = ~16'b0;
    assign data[4001] = ~16'b0;
    assign data[4002] = ~16'b0;
    assign data[4003] = ~16'b0;
    assign data[4004] = ~16'b0;
    assign data[4005] = ~16'b0;
    assign data[4006] = ~16'b0;
    assign data[4007] = ~16'b0;
    assign data[4008] = ~16'b0;
    assign data[4009] = ~16'b0;
    assign data[4010] = ~16'b0;
    assign data[4011] = ~16'b0;
    assign data[4012] = ~16'b0;
    assign data[4013] = ~16'b0;
    assign data[4014] = ~16'b0;
    assign data[4015] = ~16'b0;
    assign data[4016] = ~16'b0;
    assign data[4017] = ~16'b0;
    assign data[4018] = ~16'b0;
    assign data[4019] = ~16'b0;
    assign data[4020] = ~16'b0;
    assign data[4021] = ~16'b0;
    assign data[4022] = ~16'b0;
    assign data[4023] = ~16'b0;
    assign data[4024] = ~16'b0;
    assign data[4025] = ~16'b0;
    assign data[4026] = ~16'b0;
    assign data[4027] = ~16'b0;
    assign data[4028] = ~16'b0;
    assign data[4029] = ~16'b0;
    assign data[4030] = ~16'b0;
    assign data[4031] = ~16'b0;
    assign data[4032] = ~16'b0;
    assign data[4033] = ~16'b0;
    assign data[4034] = ~16'b0;
    assign data[4035] = ~16'b0;
    assign data[4036] = ~16'b0;
    assign data[4037] = ~16'b0;
    assign data[4038] = ~16'b0;
    assign data[4039] = ~16'b0;
    assign data[4040] = ~16'b0;
    assign data[4041] = ~16'b0;
    assign data[4042] = ~16'b0;
    assign data[4043] = ~16'b0;
    assign data[4044] = ~16'b0;
    assign data[4045] = ~16'b0;
    assign data[4046] = ~16'b0;
    assign data[4047] = ~16'b0;
    assign data[4048] = ~16'b0;
    assign data[4049] = ~16'b0;
    assign data[4050] = ~16'b0;
    assign data[4051] = ~16'b0;
    assign data[4052] = ~16'b0;
    assign data[4053] = ~16'b0;
    assign data[4054] = ~16'b0;
    assign data[4055] = ~16'b0;
    assign data[4056] = ~16'b0;
    assign data[4057] = ~16'b0;
    assign data[4058] = ~16'b0;
    assign data[4059] = ~16'b0;
    assign data[4060] = ~16'b0;
    assign data[4061] = ~16'b0;
    assign data[4062] = ~16'b0;
    assign data[4063] = ~16'b0;
    assign data[4064] = ~16'b0;
    assign data[4065] = ~16'b0;
    assign data[4066] = ~16'b0;
    assign data[4067] = ~16'b0;
    assign data[4068] = ~16'b0;
    assign data[4069] = ~16'b0;
    assign data[4070] = ~16'b0;
    assign data[4071] = ~16'b0;
    assign data[4072] = ~16'b0;
    assign data[4073] = ~16'b0;
    assign data[4074] = ~16'b0;
    assign data[4075] = ~16'b0;
    assign data[4076] = ~16'b0;
    assign data[4077] = ~16'b0;
    assign data[4078] = ~16'b0;
    assign data[4079] = ~16'b0;
    assign data[4080] = ~16'b0;
    assign data[4081] = ~16'b0;
    assign data[4082] = ~16'b0;
    assign data[4083] = ~16'b0;
    assign data[4084] = ~16'b0;
    assign data[4085] = ~16'b0;
    assign data[4086] = ~16'b0;
    assign data[4087] = ~16'b0;
    assign data[4088] = ~16'b0;
    assign data[4089] = ~16'b0;
    assign data[4090] = ~16'b0;
    assign data[4091] = ~16'b0;
    assign data[4092] = ~16'b0;
    assign data[4093] = ~16'b0;
    assign data[4094] = ~16'b0;
    assign data[4095] = ~16'b0;
    assign data[4096] = ~16'b0;
    assign data[4097] = ~16'b0;
    assign data[4098] = ~16'b0;
    assign data[4099] = ~16'b0;
    assign data[4100] = 16'b0;
    assign data[4101] = 16'b0;
    assign data[4102] = 16'b0;
    assign data[4103] = 16'b0;
    assign data[4104] = 16'b0;
    assign data[4105] = 16'b0;
    assign data[4106] = 16'b0;
    assign data[4107] = 16'b0;
    assign data[4108] = 16'b0;
    assign data[4109] = 16'b0;
    assign data[4110] = 16'b0;
    assign data[4111] = 16'b0;
    assign data[4112] = 16'b0;
    assign data[4113] = 16'b0;
    assign data[4114] = 16'b0;
    assign data[4115] = 16'b0;
    assign data[4116] = 16'b0;
    assign data[4117] = 16'b0;
    assign data[4118] = 16'b0;
    assign data[4119] = 16'b0;
    assign data[4120] = 16'b0;
    assign data[4121] = 16'b0;
    assign data[4122] = ~16'b0;
    assign data[4123] = ~16'b0;
    assign data[4124] = ~16'b0;
    assign data[4125] = ~16'b0;
    assign data[4126] = ~16'b0;
    assign data[4127] = ~16'b0;
    assign data[4128] = ~16'b0;
    assign data[4129] = ~16'b0;
    assign data[4130] = 16'b0;
    assign data[4131] = 16'b0;
    assign data[4132] = ~16'b0;
    assign data[4133] = ~16'b0;
    assign data[4134] = ~16'b0;
    assign data[4135] = ~16'b0;
    assign data[4136] = ~16'b0;
    assign data[4137] = ~16'b0;
    assign data[4138] = ~16'b0;
    assign data[4139] = ~16'b0;
    assign data[4140] = 16'b0;
    assign data[4141] = 16'b0;
    assign data[4142] = ~16'b0;
    assign data[4143] = ~16'b0;
    assign data[4144] = ~16'b0;
    assign data[4145] = ~16'b0;
    assign data[4146] = ~16'b0;
    assign data[4147] = ~16'b0;
    assign data[4148] = ~16'b0;
    assign data[4149] = ~16'b0;
    assign data[4150] = 16'b0;
    assign data[4151] = 16'b0;
    assign data[4152] = ~16'b0;
    assign data[4153] = ~16'b0;
    assign data[4154] = ~16'b0;
    assign data[4155] = ~16'b0;
    assign data[4156] = ~16'b0;
    assign data[4157] = ~16'b0;
    assign data[4158] = ~16'b0;
    assign data[4159] = ~16'b0;
    assign data[4160] = 16'b0;
    assign data[4161] = 16'b0;
    assign data[4162] = ~16'b0;
    assign data[4163] = ~16'b0;
    assign data[4164] = ~16'b0;
    assign data[4165] = ~16'b0;
    assign data[4166] = ~16'b0;
    assign data[4167] = ~16'b0;
    assign data[4168] = ~16'b0;
    assign data[4169] = ~16'b0;
    assign data[4170] = 16'b0;
    assign data[4171] = 16'b0;
    assign data[4172] = ~16'b0;
    assign data[4173] = ~16'b0;
    assign data[4174] = ~16'b0;
    assign data[4175] = ~16'b0;
    assign data[4176] = ~16'b0;
    assign data[4177] = ~16'b0;
    assign data[4178] = ~16'b0;
    assign data[4179] = ~16'b0;
    assign data[4180] = 16'b0;
    assign data[4181] = 16'b0;
    assign data[4182] = ~16'b0;
    assign data[4183] = ~16'b0;
    assign data[4184] = ~16'b0;
    assign data[4185] = ~16'b0;
    assign data[4186] = ~16'b0;
    assign data[4187] = ~16'b0;
    assign data[4188] = ~16'b0;
    assign data[4189] = ~16'b0;
    assign data[4190] = 16'b0;
    assign data[4191] = 16'b0;
    assign data[4192] = ~16'b0;
    assign data[4193] = ~16'b0;
    assign data[4194] = ~16'b0;
    assign data[4195] = ~16'b0;
    assign data[4196] = ~16'b0;
    assign data[4197] = ~16'b0;
    assign data[4198] = ~16'b0;
    assign data[4199] = ~16'b0;
    assign data[4200] = 16'b0;
    assign data[4201] = 16'b0;
    assign data[4202] = ~16'b0;
    assign data[4203] = ~16'b0;
    assign data[4204] = ~16'b0;
    assign data[4205] = ~16'b0;
    assign data[4206] = ~16'b0;
    assign data[4207] = ~16'b0;
    assign data[4208] = ~16'b0;
    assign data[4209] = ~16'b0;
    assign data[4210] = 16'b0;
    assign data[4211] = 16'b0;
    assign data[4212] = ~16'b0;
    assign data[4213] = ~16'b0;
    assign data[4214] = ~16'b0;
    assign data[4215] = ~16'b0;
    assign data[4216] = ~16'b0;
    assign data[4217] = ~16'b0;
    assign data[4218] = ~16'b0;
    assign data[4219] = ~16'b0;
    assign data[4220] = 16'b0;
    assign data[4221] = 16'b0;
    assign data[4222] = ~16'b0;
    assign data[4223] = ~16'b0;
    assign data[4224] = ~16'b0;
    assign data[4225] = ~16'b0;
    assign data[4226] = ~16'b0;
    assign data[4227] = ~16'b0;
    assign data[4228] = ~16'b0;
    assign data[4229] = ~16'b0;
    assign data[4230] = 16'b0;
    assign data[4231] = 16'b0;
    assign data[4232] = ~16'b0;
    assign data[4233] = ~16'b0;
    assign data[4234] = ~16'b0;
    assign data[4235] = ~16'b0;
    assign data[4236] = ~16'b0;
    assign data[4237] = ~16'b0;
    assign data[4238] = ~16'b0;
    assign data[4239] = ~16'b0;
    assign data[4240] = 16'b0;
    assign data[4241] = 16'b0;
    assign data[4242] = ~16'b0;
    assign data[4243] = ~16'b0;
    assign data[4244] = ~16'b0;
    assign data[4245] = ~16'b0;
    assign data[4246] = ~16'b0;
    assign data[4247] = ~16'b0;
    assign data[4248] = ~16'b0;
    assign data[4249] = ~16'b0;
    assign data[4250] = 16'b0;
    assign data[4251] = 16'b0;
    assign data[4252] = ~16'b0;
    assign data[4253] = ~16'b0;
    assign data[4254] = ~16'b0;
    assign data[4255] = ~16'b0;
    assign data[4256] = ~16'b0;
    assign data[4257] = ~16'b0;
    assign data[4258] = ~16'b0;
    assign data[4259] = ~16'b0;
    assign data[4260] = 16'b0;
    assign data[4261] = 16'b0;
    assign data[4262] = ~16'b0;
    assign data[4263] = ~16'b0;
    assign data[4264] = ~16'b0;
    assign data[4265] = ~16'b0;
    assign data[4266] = ~16'b0;
    assign data[4267] = ~16'b0;
    assign data[4268] = ~16'b0;
    assign data[4269] = ~16'b0;
    assign data[4270] = 16'b0;
    assign data[4271] = 16'b0;
    assign data[4272] = ~16'b0;
    assign data[4273] = ~16'b0;
    assign data[4274] = ~16'b0;
    assign data[4275] = ~16'b0;
    assign data[4276] = ~16'b0;
    assign data[4277] = ~16'b0;
    assign data[4278] = ~16'b0;
    assign data[4279] = ~16'b0;
    assign data[4280] = 16'b0;
    assign data[4281] = 16'b0;
    assign data[4282] = ~16'b0;
    assign data[4283] = ~16'b0;
    assign data[4284] = ~16'b0;
    assign data[4285] = ~16'b0;
    assign data[4286] = ~16'b0;
    assign data[4287] = ~16'b0;
    assign data[4288] = ~16'b0;
    assign data[4289] = ~16'b0;
    assign data[4290] = 16'b0;
    assign data[4291] = 16'b0;
    assign data[4292] = ~16'b0;
    assign data[4293] = ~16'b0;
    assign data[4294] = ~16'b0;
    assign data[4295] = ~16'b0;
    assign data[4296] = ~16'b0;
    assign data[4297] = ~16'b0;
    assign data[4298] = ~16'b0;
    assign data[4299] = ~16'b0;
    assign data[4300] = 16'b0;
    assign data[4301] = 16'b0;
    assign data[4302] = ~16'b0;
    assign data[4303] = ~16'b0;
    assign data[4304] = ~16'b0;
    assign data[4305] = ~16'b0;
    assign data[4306] = ~16'b0;
    assign data[4307] = ~16'b0;
    assign data[4308] = ~16'b0;
    assign data[4309] = ~16'b0;
    assign data[4310] = 16'b0;
    assign data[4311] = 16'b0;
    assign data[4312] = ~16'b0;
    assign data[4313] = ~16'b0;
    assign data[4314] = ~16'b0;
    assign data[4315] = ~16'b0;
    assign data[4316] = ~16'b0;
    assign data[4317] = ~16'b0;
    assign data[4318] = ~16'b0;
    assign data[4319] = ~16'b0;
    assign data[4320] = 16'b0;
    assign data[4321] = 16'b0;
    assign data[4322] = ~16'b0;
    assign data[4323] = ~16'b0;
    assign data[4324] = ~16'b0;
    assign data[4325] = ~16'b0;
    assign data[4326] = ~16'b0;
    assign data[4327] = ~16'b0;
    assign data[4328] = ~16'b0;
    assign data[4329] = ~16'b0;
    assign data[4330] = 16'b0;
    assign data[4331] = 16'b0;
    assign data[4332] = ~16'b0;
    assign data[4333] = ~16'b0;
    assign data[4334] = ~16'b0;
    assign data[4335] = ~16'b0;
    assign data[4336] = ~16'b0;
    assign data[4337] = ~16'b0;
    assign data[4338] = ~16'b0;
    assign data[4339] = ~16'b0;
    assign data[4340] = 16'b0;
    assign data[4341] = 16'b0;
    assign data[4342] = ~16'b0;
    assign data[4343] = ~16'b0;
    assign data[4344] = ~16'b0;
    assign data[4345] = ~16'b0;
    assign data[4346] = ~16'b0;
    assign data[4347] = ~16'b0;
    assign data[4348] = ~16'b0;
    assign data[4349] = ~16'b0;
    assign data[4350] = 16'b0;
    assign data[4351] = 16'b0;
    assign data[4352] = ~16'b0;
    assign data[4353] = ~16'b0;
    assign data[4354] = ~16'b0;
    assign data[4355] = ~16'b0;
    assign data[4356] = ~16'b0;
    assign data[4357] = ~16'b0;
    assign data[4358] = ~16'b0;
    assign data[4359] = ~16'b0;
    assign data[4360] = 16'b0;
    assign data[4361] = 16'b0;
    assign data[4362] = ~16'b0;
    assign data[4363] = ~16'b0;
    assign data[4364] = ~16'b0;
    assign data[4365] = ~16'b0;
    assign data[4366] = ~16'b0;
    assign data[4367] = ~16'b0;
    assign data[4368] = ~16'b0;
    assign data[4369] = ~16'b0;
    assign data[4370] = 16'b0;
    assign data[4371] = 16'b0;
    assign data[4372] = ~16'b0;
    assign data[4373] = ~16'b0;
    assign data[4374] = ~16'b0;
    assign data[4375] = ~16'b0;
    assign data[4376] = ~16'b0;
    assign data[4377] = ~16'b0;
    assign data[4378] = ~16'b0;
    assign data[4379] = ~16'b0;
    assign data[4380] = 16'b0;
    assign data[4381] = 16'b0;
    assign data[4382] = ~16'b0;
    assign data[4383] = ~16'b0;
    assign data[4384] = ~16'b0;
    assign data[4385] = ~16'b0;
    assign data[4386] = ~16'b0;
    assign data[4387] = ~16'b0;
    assign data[4388] = ~16'b0;
    assign data[4389] = ~16'b0;
    assign data[4390] = 16'b0;
    assign data[4391] = 16'b0;
    assign data[4392] = ~16'b0;
    assign data[4393] = ~16'b0;
    assign data[4394] = ~16'b0;
    assign data[4395] = ~16'b0;
    assign data[4396] = ~16'b0;
    assign data[4397] = ~16'b0;
    assign data[4398] = ~16'b0;
    assign data[4399] = ~16'b0;
    assign data[4400] = 16'b0;
    assign data[4401] = 16'b0;
    assign data[4402] = ~16'b0;
    assign data[4403] = ~16'b0;
    assign data[4404] = ~16'b0;
    assign data[4405] = ~16'b0;
    assign data[4406] = ~16'b0;
    assign data[4407] = ~16'b0;
    assign data[4408] = ~16'b0;
    assign data[4409] = ~16'b0;
    assign data[4410] = 16'b0;
    assign data[4411] = 16'b0;
    assign data[4412] = ~16'b0;
    assign data[4413] = ~16'b0;
    assign data[4414] = ~16'b0;
    assign data[4415] = ~16'b0;
    assign data[4416] = ~16'b0;
    assign data[4417] = ~16'b0;
    assign data[4418] = ~16'b0;
    assign data[4419] = ~16'b0;
    assign data[4420] = 16'b0;
    assign data[4421] = 16'b0;
    assign data[4422] = ~16'b0;
    assign data[4423] = ~16'b0;
    assign data[4424] = ~16'b0;
    assign data[4425] = ~16'b0;
    assign data[4426] = ~16'b0;
    assign data[4427] = ~16'b0;
    assign data[4428] = ~16'b0;
    assign data[4429] = ~16'b0;
    assign data[4430] = 16'b0;
    assign data[4431] = 16'b0;
    assign data[4432] = ~16'b0;
    assign data[4433] = ~16'b0;
    assign data[4434] = ~16'b0;
    assign data[4435] = ~16'b0;
    assign data[4436] = ~16'b0;
    assign data[4437] = ~16'b0;
    assign data[4438] = ~16'b0;
    assign data[4439] = ~16'b0;
    assign data[4440] = 16'b0;
    assign data[4441] = 16'b0;
    assign data[4442] = 16'b0;
    assign data[4443] = 16'b0;
    assign data[4444] = 16'b0;
    assign data[4445] = 16'b0;
    assign data[4446] = 16'b0;
    assign data[4447] = 16'b0;
    assign data[4448] = 16'b0;
    assign data[4449] = 16'b0;
    assign data[4450] = 16'b0;
    assign data[4451] = 16'b0;
    assign data[4452] = 16'b0;
    assign data[4453] = 16'b0;
    assign data[4454] = 16'b0;
    assign data[4455] = 16'b0;
    assign data[4456] = 16'b0;
    assign data[4457] = 16'b0;
    assign data[4458] = 16'b0;
    assign data[4459] = 16'b0;
    assign data[4460] = ~16'b0;
    assign data[4461] = ~16'b0;
    assign data[4462] = ~16'b0;
    assign data[4463] = ~16'b0;
    assign data[4464] = ~16'b0;
    assign data[4465] = ~16'b0;
    assign data[4466] = ~16'b0;
    assign data[4467] = ~16'b0;
    assign data[4468] = ~16'b0;
    assign data[4469] = ~16'b0;
    assign data[4470] = ~16'b0;
    assign data[4471] = ~16'b0;
    assign data[4472] = ~16'b0;
    assign data[4473] = ~16'b0;
    assign data[4474] = ~16'b0;
    assign data[4475] = ~16'b0;
    assign data[4476] = ~16'b0;
    assign data[4477] = ~16'b0;
    assign data[4478] = ~16'b0;
    assign data[4479] = ~16'b0;
    assign data[4480] = ~16'b0;
    assign data[4481] = ~16'b0;
    assign data[4482] = ~16'b0;
    assign data[4483] = ~16'b0;
    assign data[4484] = ~16'b0;
    assign data[4485] = ~16'b0;
    assign data[4486] = ~16'b0;
    assign data[4487] = ~16'b0;
    assign data[4488] = ~16'b0;
    assign data[4489] = ~16'b0;
    assign data[4490] = ~16'b0;
    assign data[4491] = ~16'b0;
    assign data[4492] = ~16'b0;
    assign data[4493] = ~16'b0;
    assign data[4494] = ~16'b0;
    assign data[4495] = ~16'b0;
    assign data[4496] = ~16'b0;
    assign data[4497] = ~16'b0;
    assign data[4498] = ~16'b0;
    assign data[4499] = ~16'b0;
    assign data[4500] = ~16'b0;
    assign data[4501] = ~16'b0;
    assign data[4502] = ~16'b0;
    assign data[4503] = ~16'b0;
    assign data[4504] = ~16'b0;
    assign data[4505] = ~16'b0;
    assign data[4506] = ~16'b0;
    assign data[4507] = ~16'b0;
    assign data[4508] = ~16'b0;
    assign data[4509] = ~16'b0;
    assign data[4510] = ~16'b0;
    assign data[4511] = ~16'b0;
    assign data[4512] = ~16'b0;
    assign data[4513] = ~16'b0;
    assign data[4514] = ~16'b0;
    assign data[4515] = ~16'b0;
    assign data[4516] = ~16'b0;
    assign data[4517] = ~16'b0;
    assign data[4518] = ~16'b0;
    assign data[4519] = ~16'b0;
    assign data[4520] = ~16'b0;
    assign data[4521] = ~16'b0;
    assign data[4522] = ~16'b0;
    assign data[4523] = ~16'b0;
    assign data[4524] = ~16'b0;
    assign data[4525] = ~16'b0;
    assign data[4526] = ~16'b0;
    assign data[4527] = ~16'b0;
    assign data[4528] = ~16'b0;
    assign data[4529] = ~16'b0;
    assign data[4530] = ~16'b0;
    assign data[4531] = ~16'b0;
    assign data[4532] = ~16'b0;
    assign data[4533] = ~16'b0;
    assign data[4534] = ~16'b0;
    assign data[4535] = ~16'b0;
    assign data[4536] = ~16'b0;
    assign data[4537] = ~16'b0;
    assign data[4538] = ~16'b0;
    assign data[4539] = ~16'b0;
    assign data[4540] = ~16'b0;
    assign data[4541] = ~16'b0;
    assign data[4542] = ~16'b0;
    assign data[4543] = ~16'b0;
    assign data[4544] = ~16'b0;
    assign data[4545] = ~16'b0;
    assign data[4546] = ~16'b0;
    assign data[4547] = ~16'b0;
    assign data[4548] = ~16'b0;
    assign data[4549] = ~16'b0;
    assign data[4550] = ~16'b0;
    assign data[4551] = ~16'b0;
    assign data[4552] = ~16'b0;
    assign data[4553] = ~16'b0;
    assign data[4554] = ~16'b0;
    assign data[4555] = ~16'b0;
    assign data[4556] = ~16'b0;
    assign data[4557] = ~16'b0;
    assign data[4558] = ~16'b0;
    assign data[4559] = ~16'b0;
    assign data[4560] = ~16'b0;
    assign data[4561] = ~16'b0;
    assign data[4562] = ~16'b0;
    assign data[4563] = ~16'b0;
    assign data[4564] = ~16'b0;
    assign data[4565] = ~16'b0;
    assign data[4566] = ~16'b0;
    assign data[4567] = ~16'b0;
    assign data[4568] = ~16'b0;
    assign data[4569] = ~16'b0;
    assign data[4570] = ~16'b0;
    assign data[4571] = ~16'b0;
    assign data[4572] = ~16'b0;
    assign data[4573] = ~16'b0;
    assign data[4574] = ~16'b0;
    assign data[4575] = ~16'b0;
    assign data[4576] = ~16'b0;
    assign data[4577] = ~16'b0;
    assign data[4578] = ~16'b0;
    assign data[4579] = ~16'b0;
    assign data[4580] = ~16'b0;
    assign data[4581] = ~16'b0;
    assign data[4582] = ~16'b0;
    assign data[4583] = ~16'b0;
    assign data[4584] = ~16'b0;
    assign data[4585] = ~16'b0;
    assign data[4586] = ~16'b0;
    assign data[4587] = ~16'b0;
    assign data[4588] = ~16'b0;
    assign data[4589] = ~16'b0;
    assign data[4590] = ~16'b0;
    assign data[4591] = ~16'b0;
    assign data[4592] = ~16'b0;
    assign data[4593] = ~16'b0;
    assign data[4594] = ~16'b0;
    assign data[4595] = ~16'b0;
    assign data[4596] = ~16'b0;
    assign data[4597] = ~16'b0;
    assign data[4598] = ~16'b0;
    assign data[4599] = ~16'b0;
    assign data[4600] = ~16'b0;
    assign data[4601] = ~16'b0;
    assign data[4602] = ~16'b0;
    assign data[4603] = ~16'b0;
    assign data[4604] = ~16'b0;
    assign data[4605] = ~16'b0;
    assign data[4606] = ~16'b0;
    assign data[4607] = ~16'b0;
    assign data[4608] = ~16'b0;
    assign data[4609] = ~16'b0;
    assign data[4610] = ~16'b0;
    assign data[4611] = ~16'b0;
    assign data[4612] = ~16'b0;
    assign data[4613] = ~16'b0;
    assign data[4614] = ~16'b0;
    assign data[4615] = ~16'b0;
    assign data[4616] = ~16'b0;
    assign data[4617] = ~16'b0;
    assign data[4618] = ~16'b0;
    assign data[4619] = ~16'b0;
    assign data[4620] = ~16'b0;
    assign data[4621] = ~16'b0;
    assign data[4622] = ~16'b0;
    assign data[4623] = ~16'b0;
    assign data[4624] = ~16'b0;
    assign data[4625] = ~16'b0;
    assign data[4626] = ~16'b0;
    assign data[4627] = ~16'b0;
    assign data[4628] = ~16'b0;
    assign data[4629] = ~16'b0;
    assign data[4630] = ~16'b0;
    assign data[4631] = ~16'b0;
    assign data[4632] = ~16'b0;
    assign data[4633] = ~16'b0;
    assign data[4634] = ~16'b0;
    assign data[4635] = ~16'b0;
    assign data[4636] = ~16'b0;
    assign data[4637] = ~16'b0;
    assign data[4638] = ~16'b0;
    assign data[4639] = ~16'b0;
    assign data[4640] = ~16'b0;
    assign data[4641] = ~16'b0;
    assign data[4642] = ~16'b0;
    assign data[4643] = ~16'b0;
    assign data[4644] = ~16'b0;
    assign data[4645] = ~16'b0;
    assign data[4646] = ~16'b0;
    assign data[4647] = ~16'b0;
    assign data[4648] = ~16'b0;
    assign data[4649] = ~16'b0;
    assign data[4650] = ~16'b0;
    assign data[4651] = ~16'b0;
    assign data[4652] = ~16'b0;
    assign data[4653] = ~16'b0;
    assign data[4654] = ~16'b0;
    assign data[4655] = ~16'b0;
    assign data[4656] = ~16'b0;
    assign data[4657] = ~16'b0;
    assign data[4658] = ~16'b0;
    assign data[4659] = ~16'b0;
    assign data[4660] = ~16'b0;
    assign data[4661] = ~16'b0;
    assign data[4662] = ~16'b0;
    assign data[4663] = ~16'b0;
    assign data[4664] = ~16'b0;
    assign data[4665] = ~16'b0;
    assign data[4666] = ~16'b0;
    assign data[4667] = ~16'b0;
    assign data[4668] = ~16'b0;
    assign data[4669] = ~16'b0;
    assign data[4670] = ~16'b0;
    assign data[4671] = ~16'b0;
    assign data[4672] = ~16'b0;
    assign data[4673] = ~16'b0;
    assign data[4674] = ~16'b0;
    assign data[4675] = ~16'b0;
    assign data[4676] = ~16'b0;
    assign data[4677] = ~16'b0;
    assign data[4678] = ~16'b0;
    assign data[4679] = ~16'b0;
    assign data[4680] = ~16'b0;
    assign data[4681] = ~16'b0;
    assign data[4682] = ~16'b0;
    assign data[4683] = ~16'b0;
    assign data[4684] = ~16'b0;
    assign data[4685] = ~16'b0;
    assign data[4686] = ~16'b0;
    assign data[4687] = ~16'b0;
    assign data[4688] = ~16'b0;
    assign data[4689] = ~16'b0;
    assign data[4690] = ~16'b0;
    assign data[4691] = ~16'b0;
    assign data[4692] = ~16'b0;
    assign data[4693] = ~16'b0;
    assign data[4694] = ~16'b0;
    assign data[4695] = ~16'b0;
    assign data[4696] = ~16'b0;
    assign data[4697] = ~16'b0;
    assign data[4698] = ~16'b0;
    assign data[4699] = ~16'b0;
    assign data[4700] = ~16'b0;
    assign data[4701] = ~16'b0;
    assign data[4702] = ~16'b0;
    assign data[4703] = ~16'b0;
    assign data[4704] = ~16'b0;
    assign data[4705] = ~16'b0;
    assign data[4706] = ~16'b0;
    assign data[4707] = ~16'b0;
    assign data[4708] = ~16'b0;
    assign data[4709] = ~16'b0;
    assign data[4710] = ~16'b0;
    assign data[4711] = ~16'b0;
    assign data[4712] = ~16'b0;
    assign data[4713] = ~16'b0;
    assign data[4714] = ~16'b0;
    assign data[4715] = ~16'b0;
    assign data[4716] = ~16'b0;
    assign data[4717] = ~16'b0;
    assign data[4718] = ~16'b0;
    assign data[4719] = ~16'b0;
    assign data[4720] = ~16'b0;
    assign data[4721] = ~16'b0;
    assign data[4722] = ~16'b0;
    assign data[4723] = ~16'b0;
    assign data[4724] = ~16'b0;
    assign data[4725] = ~16'b0;
    assign data[4726] = ~16'b0;
    assign data[4727] = ~16'b0;
    assign data[4728] = ~16'b0;
    assign data[4729] = ~16'b0;
    assign data[4730] = ~16'b0;
    assign data[4731] = ~16'b0;
    assign data[4732] = ~16'b0;
    assign data[4733] = ~16'b0;
    assign data[4734] = ~16'b0;
    assign data[4735] = ~16'b0;
    assign data[4736] = ~16'b0;
    assign data[4737] = ~16'b0;
    assign data[4738] = ~16'b0;
    assign data[4739] = ~16'b0;
    assign data[4740] = ~16'b0;
    assign data[4741] = ~16'b0;
    assign data[4742] = ~16'b0;
    assign data[4743] = ~16'b0;
    assign data[4744] = ~16'b0;
    assign data[4745] = ~16'b0;
    assign data[4746] = ~16'b0;
    assign data[4747] = ~16'b0;
    assign data[4748] = ~16'b0;
    assign data[4749] = ~16'b0;
    assign data[4750] = ~16'b0;
    assign data[4751] = ~16'b0;
    assign data[4752] = ~16'b0;
    assign data[4753] = ~16'b0;
    assign data[4754] = ~16'b0;
    assign data[4755] = ~16'b0;
    assign data[4756] = ~16'b0;
    assign data[4757] = ~16'b0;
    assign data[4758] = ~16'b0;
    assign data[4759] = ~16'b0;
    assign data[4760] = ~16'b0;
    assign data[4761] = ~16'b0;
    assign data[4762] = ~16'b0;
    assign data[4763] = ~16'b0;
    assign data[4764] = ~16'b0;
    assign data[4765] = ~16'b0;
    assign data[4766] = ~16'b0;
    assign data[4767] = ~16'b0;
    assign data[4768] = ~16'b0;
    assign data[4769] = ~16'b0;
    assign data[4770] = ~16'b0;
    assign data[4771] = ~16'b0;
    assign data[4772] = ~16'b0;
    assign data[4773] = ~16'b0;
    assign data[4774] = ~16'b0;
    assign data[4775] = ~16'b0;
    assign data[4776] = ~16'b0;
    assign data[4777] = ~16'b0;
    assign data[4778] = ~16'b0;
    assign data[4779] = ~16'b0;
    assign data[4780] = ~16'b0;
    assign data[4781] = ~16'b0;
    assign data[4782] = ~16'b0;
    assign data[4783] = ~16'b0;
    assign data[4784] = ~16'b0;
    assign data[4785] = ~16'b0;
    assign data[4786] = ~16'b0;
    assign data[4787] = ~16'b0;
    assign data[4788] = ~16'b0;
    assign data[4789] = ~16'b0;
    assign data[4790] = ~16'b0;
    assign data[4791] = ~16'b0;
    assign data[4792] = ~16'b0;
    assign data[4793] = ~16'b0;
    assign data[4794] = ~16'b0;
    assign data[4795] = ~16'b0;
    assign data[4796] = ~16'b0;
    assign data[4797] = ~16'b0;
    assign data[4798] = ~16'b0;
    assign data[4799] = ~16'b0;
    assign data[4800] = ~16'b0;
    assign data[4801] = ~16'b0;
    assign data[4802] = ~16'b0;
    assign data[4803] = ~16'b0;
    assign data[4804] = ~16'b0;
    assign data[4805] = ~16'b0;
    assign data[4806] = ~16'b0;
    assign data[4807] = ~16'b0;
    assign data[4808] = ~16'b0;
    assign data[4809] = ~16'b0;
    assign data[4810] = ~16'b0;
    assign data[4811] = ~16'b0;
    assign data[4812] = ~16'b0;
    assign data[4813] = ~16'b0;
    assign data[4814] = ~16'b0;
    assign data[4815] = ~16'b0;
    assign data[4816] = ~16'b0;
    assign data[4817] = ~16'b0;
    assign data[4818] = ~16'b0;
    assign data[4819] = ~16'b0;
    assign data[4820] = 16'b0;
    assign data[4821] = 16'b0;
    assign data[4822] = 16'b0;
    assign data[4823] = 16'b0;
    assign data[4824] = 16'b0;
    assign data[4825] = 16'b0;
    assign data[4826] = 16'b0;
    assign data[4827] = 16'b0;
    assign data[4828] = 16'b0;
    assign data[4829] = 16'b0;
    assign data[4830] = 16'b0;
    assign data[4831] = 16'b0;
    assign data[4832] = 16'b0;
    assign data[4833] = 16'b0;
    assign data[4834] = 16'b0;
    assign data[4835] = 16'b0;
    assign data[4836] = 16'b0;
    assign data[4837] = 16'b0;
    assign data[4838] = 16'b0;
    assign data[4839] = 16'b0;
    assign data[4840] = 16'b0;
    assign data[4841] = 16'b0;
    assign data[4842] = ~16'b0;
    assign data[4843] = ~16'b0;
    assign data[4844] = ~16'b0;
    assign data[4845] = ~16'b0;
    assign data[4846] = ~16'b0;
    assign data[4847] = ~16'b0;
    assign data[4848] = ~16'b0;
    assign data[4849] = ~16'b0;
    assign data[4850] = 16'b0;
    assign data[4851] = 16'b0;
    assign data[4852] = ~16'b0;
    assign data[4853] = ~16'b0;
    assign data[4854] = ~16'b0;
    assign data[4855] = ~16'b0;
    assign data[4856] = ~16'b0;
    assign data[4857] = ~16'b0;
    assign data[4858] = ~16'b0;
    assign data[4859] = ~16'b0;
    assign data[4860] = 16'b0;
    assign data[4861] = 16'b0;
    assign data[4862] = ~16'b0;
    assign data[4863] = ~16'b0;
    assign data[4864] = ~16'b0;
    assign data[4865] = ~16'b0;
    assign data[4866] = ~16'b0;
    assign data[4867] = ~16'b0;
    assign data[4868] = ~16'b0;
    assign data[4869] = ~16'b0;
    assign data[4870] = 16'b0;
    assign data[4871] = 16'b0;
    assign data[4872] = ~16'b0;
    assign data[4873] = ~16'b0;
    assign data[4874] = ~16'b0;
    assign data[4875] = ~16'b0;
    assign data[4876] = ~16'b0;
    assign data[4877] = ~16'b0;
    assign data[4878] = ~16'b0;
    assign data[4879] = ~16'b0;
    assign data[4880] = 16'b0;
    assign data[4881] = 16'b0;
    assign data[4882] = ~16'b0;
    assign data[4883] = ~16'b0;
    assign data[4884] = ~16'b0;
    assign data[4885] = ~16'b0;
    assign data[4886] = ~16'b0;
    assign data[4887] = ~16'b0;
    assign data[4888] = ~16'b0;
    assign data[4889] = ~16'b0;
    assign data[4890] = 16'b0;
    assign data[4891] = 16'b0;
    assign data[4892] = ~16'b0;
    assign data[4893] = ~16'b0;
    assign data[4894] = ~16'b0;
    assign data[4895] = ~16'b0;
    assign data[4896] = ~16'b0;
    assign data[4897] = ~16'b0;
    assign data[4898] = ~16'b0;
    assign data[4899] = ~16'b0;
    assign data[4900] = 16'b0;
    assign data[4901] = 16'b0;
    assign data[4902] = ~16'b0;
    assign data[4903] = ~16'b0;
    assign data[4904] = ~16'b0;
    assign data[4905] = ~16'b0;
    assign data[4906] = ~16'b0;
    assign data[4907] = ~16'b0;
    assign data[4908] = ~16'b0;
    assign data[4909] = ~16'b0;
    assign data[4910] = 16'b0;
    assign data[4911] = 16'b0;
    assign data[4912] = ~16'b0;
    assign data[4913] = ~16'b0;
    assign data[4914] = ~16'b0;
    assign data[4915] = ~16'b0;
    assign data[4916] = ~16'b0;
    assign data[4917] = ~16'b0;
    assign data[4918] = ~16'b0;
    assign data[4919] = ~16'b0;
    assign data[4920] = 16'b0;
    assign data[4921] = 16'b0;
    assign data[4922] = ~16'b0;
    assign data[4923] = ~16'b0;
    assign data[4924] = ~16'b0;
    assign data[4925] = ~16'b0;
    assign data[4926] = ~16'b0;
    assign data[4927] = ~16'b0;
    assign data[4928] = ~16'b0;
    assign data[4929] = ~16'b0;
    assign data[4930] = 16'b0;
    assign data[4931] = 16'b0;
    assign data[4932] = ~16'b0;
    assign data[4933] = ~16'b0;
    assign data[4934] = ~16'b0;
    assign data[4935] = ~16'b0;
    assign data[4936] = ~16'b0;
    assign data[4937] = ~16'b0;
    assign data[4938] = ~16'b0;
    assign data[4939] = ~16'b0;
    assign data[4940] = 16'b0;
    assign data[4941] = 16'b0;
    assign data[4942] = ~16'b0;
    assign data[4943] = ~16'b0;
    assign data[4944] = ~16'b0;
    assign data[4945] = ~16'b0;
    assign data[4946] = ~16'b0;
    assign data[4947] = ~16'b0;
    assign data[4948] = ~16'b0;
    assign data[4949] = ~16'b0;
    assign data[4950] = 16'b0;
    assign data[4951] = 16'b0;
    assign data[4952] = ~16'b0;
    assign data[4953] = ~16'b0;
    assign data[4954] = ~16'b0;
    assign data[4955] = ~16'b0;
    assign data[4956] = ~16'b0;
    assign data[4957] = ~16'b0;
    assign data[4958] = ~16'b0;
    assign data[4959] = ~16'b0;
    assign data[4960] = 16'b0;
    assign data[4961] = 16'b0;
    assign data[4962] = ~16'b0;
    assign data[4963] = ~16'b0;
    assign data[4964] = ~16'b0;
    assign data[4965] = ~16'b0;
    assign data[4966] = ~16'b0;
    assign data[4967] = ~16'b0;
    assign data[4968] = ~16'b0;
    assign data[4969] = ~16'b0;
    assign data[4970] = 16'b0;
    assign data[4971] = 16'b0;
    assign data[4972] = ~16'b0;
    assign data[4973] = ~16'b0;
    assign data[4974] = ~16'b0;
    assign data[4975] = ~16'b0;
    assign data[4976] = ~16'b0;
    assign data[4977] = ~16'b0;
    assign data[4978] = ~16'b0;
    assign data[4979] = ~16'b0;
    assign data[4980] = 16'b0;
    assign data[4981] = 16'b0;
    assign data[4982] = ~16'b0;
    assign data[4983] = ~16'b0;
    assign data[4984] = ~16'b0;
    assign data[4985] = ~16'b0;
    assign data[4986] = ~16'b0;
    assign data[4987] = ~16'b0;
    assign data[4988] = ~16'b0;
    assign data[4989] = ~16'b0;
    assign data[4990] = 16'b0;
    assign data[4991] = 16'b0;
    assign data[4992] = ~16'b0;
    assign data[4993] = ~16'b0;
    assign data[4994] = ~16'b0;
    assign data[4995] = ~16'b0;
    assign data[4996] = ~16'b0;
    assign data[4997] = ~16'b0;
    assign data[4998] = ~16'b0;
    assign data[4999] = ~16'b0;
    assign data[5000] = 16'b0;
    assign data[5001] = 16'b0;
    assign data[5002] = ~16'b0;
    assign data[5003] = ~16'b0;
    assign data[5004] = ~16'b0;
    assign data[5005] = ~16'b0;
    assign data[5006] = ~16'b0;
    assign data[5007] = ~16'b0;
    assign data[5008] = ~16'b0;
    assign data[5009] = ~16'b0;
    assign data[5010] = 16'b0;
    assign data[5011] = 16'b0;
    assign data[5012] = ~16'b0;
    assign data[5013] = ~16'b0;
    assign data[5014] = ~16'b0;
    assign data[5015] = ~16'b0;
    assign data[5016] = ~16'b0;
    assign data[5017] = ~16'b0;
    assign data[5018] = ~16'b0;
    assign data[5019] = ~16'b0;
    assign data[5020] = 16'b0;
    assign data[5021] = 16'b0;
    assign data[5022] = ~16'b0;
    assign data[5023] = ~16'b0;
    assign data[5024] = ~16'b0;
    assign data[5025] = ~16'b0;
    assign data[5026] = ~16'b0;
    assign data[5027] = ~16'b0;
    assign data[5028] = ~16'b0;
    assign data[5029] = ~16'b0;
    assign data[5030] = 16'b0;
    assign data[5031] = 16'b0;
    assign data[5032] = ~16'b0;
    assign data[5033] = ~16'b0;
    assign data[5034] = ~16'b0;
    assign data[5035] = ~16'b0;
    assign data[5036] = ~16'b0;
    assign data[5037] = ~16'b0;
    assign data[5038] = ~16'b0;
    assign data[5039] = ~16'b0;
    assign data[5040] = 16'b0;
    assign data[5041] = 16'b0;
    assign data[5042] = ~16'b0;
    assign data[5043] = ~16'b0;
    assign data[5044] = ~16'b0;
    assign data[5045] = ~16'b0;
    assign data[5046] = ~16'b0;
    assign data[5047] = ~16'b0;
    assign data[5048] = ~16'b0;
    assign data[5049] = ~16'b0;
    assign data[5050] = 16'b0;
    assign data[5051] = 16'b0;
    assign data[5052] = ~16'b0;
    assign data[5053] = ~16'b0;
    assign data[5054] = ~16'b0;
    assign data[5055] = ~16'b0;
    assign data[5056] = ~16'b0;
    assign data[5057] = ~16'b0;
    assign data[5058] = ~16'b0;
    assign data[5059] = ~16'b0;
    assign data[5060] = 16'b0;
    assign data[5061] = 16'b0;
    assign data[5062] = ~16'b0;
    assign data[5063] = ~16'b0;
    assign data[5064] = ~16'b0;
    assign data[5065] = ~16'b0;
    assign data[5066] = ~16'b0;
    assign data[5067] = ~16'b0;
    assign data[5068] = ~16'b0;
    assign data[5069] = ~16'b0;
    assign data[5070] = 16'b0;
    assign data[5071] = 16'b0;
    assign data[5072] = ~16'b0;
    assign data[5073] = ~16'b0;
    assign data[5074] = ~16'b0;
    assign data[5075] = ~16'b0;
    assign data[5076] = ~16'b0;
    assign data[5077] = ~16'b0;
    assign data[5078] = ~16'b0;
    assign data[5079] = ~16'b0;
    assign data[5080] = 16'b0;
    assign data[5081] = 16'b0;
    assign data[5082] = ~16'b0;
    assign data[5083] = ~16'b0;
    assign data[5084] = ~16'b0;
    assign data[5085] = ~16'b0;
    assign data[5086] = ~16'b0;
    assign data[5087] = ~16'b0;
    assign data[5088] = ~16'b0;
    assign data[5089] = ~16'b0;
    assign data[5090] = 16'b0;
    assign data[5091] = 16'b0;
    assign data[5092] = ~16'b0;
    assign data[5093] = ~16'b0;
    assign data[5094] = ~16'b0;
    assign data[5095] = ~16'b0;
    assign data[5096] = ~16'b0;
    assign data[5097] = ~16'b0;
    assign data[5098] = ~16'b0;
    assign data[5099] = ~16'b0;
    assign data[5100] = 16'b0;
    assign data[5101] = 16'b0;
    assign data[5102] = ~16'b0;
    assign data[5103] = ~16'b0;
    assign data[5104] = ~16'b0;
    assign data[5105] = ~16'b0;
    assign data[5106] = ~16'b0;
    assign data[5107] = ~16'b0;
    assign data[5108] = ~16'b0;
    assign data[5109] = ~16'b0;
    assign data[5110] = 16'b0;
    assign data[5111] = 16'b0;
    assign data[5112] = ~16'b0;
    assign data[5113] = ~16'b0;
    assign data[5114] = ~16'b0;
    assign data[5115] = ~16'b0;
    assign data[5116] = ~16'b0;
    assign data[5117] = ~16'b0;
    assign data[5118] = ~16'b0;
    assign data[5119] = ~16'b0;
    assign data[5120] = 16'b0;
    assign data[5121] = 16'b0;
    assign data[5122] = ~16'b0;
    assign data[5123] = ~16'b0;
    assign data[5124] = ~16'b0;
    assign data[5125] = ~16'b0;
    assign data[5126] = ~16'b0;
    assign data[5127] = ~16'b0;
    assign data[5128] = ~16'b0;
    assign data[5129] = ~16'b0;
    assign data[5130] = 16'b0;
    assign data[5131] = 16'b0;
    assign data[5132] = ~16'b0;
    assign data[5133] = ~16'b0;
    assign data[5134] = ~16'b0;
    assign data[5135] = ~16'b0;
    assign data[5136] = ~16'b0;
    assign data[5137] = ~16'b0;
    assign data[5138] = ~16'b0;
    assign data[5139] = ~16'b0;
    assign data[5140] = 16'b0;
    assign data[5141] = 16'b0;
    assign data[5142] = ~16'b0;
    assign data[5143] = ~16'b0;
    assign data[5144] = ~16'b0;
    assign data[5145] = ~16'b0;
    assign data[5146] = ~16'b0;
    assign data[5147] = ~16'b0;
    assign data[5148] = ~16'b0;
    assign data[5149] = ~16'b0;
    assign data[5150] = 16'b0;
    assign data[5151] = 16'b0;
    assign data[5152] = ~16'b0;
    assign data[5153] = ~16'b0;
    assign data[5154] = ~16'b0;
    assign data[5155] = ~16'b0;
    assign data[5156] = ~16'b0;
    assign data[5157] = ~16'b0;
    assign data[5158] = ~16'b0;
    assign data[5159] = ~16'b0;
    assign data[5160] = 16'b0;
    assign data[5161] = 16'b0;
    assign data[5162] = ~16'b0;
    assign data[5163] = ~16'b0;
    assign data[5164] = ~16'b0;
    assign data[5165] = ~16'b0;
    assign data[5166] = ~16'b0;
    assign data[5167] = ~16'b0;
    assign data[5168] = ~16'b0;
    assign data[5169] = ~16'b0;
    assign data[5170] = 16'b0;
    assign data[5171] = 16'b0;
    assign data[5172] = ~16'b0;
    assign data[5173] = ~16'b0;
    assign data[5174] = ~16'b0;
    assign data[5175] = ~16'b0;
    assign data[5176] = ~16'b0;
    assign data[5177] = ~16'b0;
    assign data[5178] = ~16'b0;
    assign data[5179] = ~16'b0;
    assign data[5180] = 16'b0;
    assign data[5181] = 16'b0;
    assign data[5182] = ~16'b0;
    assign data[5183] = ~16'b0;
    assign data[5184] = ~16'b0;
    assign data[5185] = ~16'b0;
    assign data[5186] = ~16'b0;
    assign data[5187] = ~16'b0;
    assign data[5188] = ~16'b0;
    assign data[5189] = ~16'b0;
    assign data[5190] = 16'b0;
    assign data[5191] = 16'b0;
    assign data[5192] = ~16'b0;
    assign data[5193] = ~16'b0;
    assign data[5194] = ~16'b0;
    assign data[5195] = ~16'b0;
    assign data[5196] = ~16'b0;
    assign data[5197] = ~16'b0;
    assign data[5198] = ~16'b0;
    assign data[5199] = ~16'b0;
    assign data[5200] = 16'b0;
    assign data[5201] = 16'b0;
    assign data[5202] = ~16'b0;
    assign data[5203] = ~16'b0;
    assign data[5204] = ~16'b0;
    assign data[5205] = ~16'b0;
    assign data[5206] = ~16'b0;
    assign data[5207] = ~16'b0;
    assign data[5208] = ~16'b0;
    assign data[5209] = ~16'b0;
    assign data[5210] = 16'b0;
    assign data[5211] = 16'b0;
    assign data[5212] = ~16'b0;
    assign data[5213] = ~16'b0;
    assign data[5214] = ~16'b0;
    assign data[5215] = ~16'b0;
    assign data[5216] = ~16'b0;
    assign data[5217] = ~16'b0;
    assign data[5218] = ~16'b0;
    assign data[5219] = ~16'b0;
    assign data[5220] = 16'b0;
    assign data[5221] = 16'b0;
    assign data[5222] = ~16'b0;
    assign data[5223] = ~16'b0;
    assign data[5224] = ~16'b0;
    assign data[5225] = ~16'b0;
    assign data[5226] = ~16'b0;
    assign data[5227] = ~16'b0;
    assign data[5228] = ~16'b0;
    assign data[5229] = ~16'b0;
    assign data[5230] = 16'b0;
    assign data[5231] = 16'b0;
    assign data[5232] = ~16'b0;
    assign data[5233] = ~16'b0;
    assign data[5234] = ~16'b0;
    assign data[5235] = ~16'b0;
    assign data[5236] = ~16'b0;
    assign data[5237] = ~16'b0;
    assign data[5238] = ~16'b0;
    assign data[5239] = ~16'b0;
    assign data[5240] = 16'b0;
    assign data[5241] = 16'b0;
    assign data[5242] = ~16'b0;
    assign data[5243] = ~16'b0;
    assign data[5244] = ~16'b0;
    assign data[5245] = ~16'b0;
    assign data[5246] = ~16'b0;
    assign data[5247] = ~16'b0;
    assign data[5248] = ~16'b0;
    assign data[5249] = ~16'b0;
    assign data[5250] = 16'b0;
    assign data[5251] = 16'b0;
    assign data[5252] = ~16'b0;
    assign data[5253] = ~16'b0;
    assign data[5254] = ~16'b0;
    assign data[5255] = ~16'b0;
    assign data[5256] = ~16'b0;
    assign data[5257] = ~16'b0;
    assign data[5258] = ~16'b0;
    assign data[5259] = ~16'b0;
    assign data[5260] = 16'b0;
    assign data[5261] = 16'b0;
    assign data[5262] = ~16'b0;
    assign data[5263] = ~16'b0;
    assign data[5264] = ~16'b0;
    assign data[5265] = ~16'b0;
    assign data[5266] = ~16'b0;
    assign data[5267] = ~16'b0;
    assign data[5268] = ~16'b0;
    assign data[5269] = ~16'b0;
    assign data[5270] = 16'b0;
    assign data[5271] = 16'b0;
    assign data[5272] = ~16'b0;
    assign data[5273] = ~16'b0;
    assign data[5274] = ~16'b0;
    assign data[5275] = ~16'b0;
    assign data[5276] = ~16'b0;
    assign data[5277] = ~16'b0;
    assign data[5278] = ~16'b0;
    assign data[5279] = ~16'b0;
    assign data[5280] = 16'b0;
    assign data[5281] = 16'b0;
    assign data[5282] = ~16'b0;
    assign data[5283] = ~16'b0;
    assign data[5284] = ~16'b0;
    assign data[5285] = ~16'b0;
    assign data[5286] = ~16'b0;
    assign data[5287] = ~16'b0;
    assign data[5288] = ~16'b0;
    assign data[5289] = ~16'b0;
    assign data[5290] = 16'b0;
    assign data[5291] = 16'b0;
    assign data[5292] = ~16'b0;
    assign data[5293] = ~16'b0;
    assign data[5294] = ~16'b0;
    assign data[5295] = ~16'b0;
    assign data[5296] = ~16'b0;
    assign data[5297] = ~16'b0;
    assign data[5298] = ~16'b0;
    assign data[5299] = ~16'b0;
    assign data[5300] = 16'b0;
    assign data[5301] = 16'b0;
    assign data[5302] = ~16'b0;
    assign data[5303] = ~16'b0;
    assign data[5304] = ~16'b0;
    assign data[5305] = ~16'b0;
    assign data[5306] = ~16'b0;
    assign data[5307] = ~16'b0;
    assign data[5308] = ~16'b0;
    assign data[5309] = ~16'b0;
    assign data[5310] = 16'b0;
    assign data[5311] = 16'b0;
    assign data[5312] = ~16'b0;
    assign data[5313] = ~16'b0;
    assign data[5314] = ~16'b0;
    assign data[5315] = ~16'b0;
    assign data[5316] = ~16'b0;
    assign data[5317] = ~16'b0;
    assign data[5318] = ~16'b0;
    assign data[5319] = ~16'b0;
    assign data[5320] = 16'b0;
    assign data[5321] = 16'b0;
    assign data[5322] = ~16'b0;
    assign data[5323] = ~16'b0;
    assign data[5324] = ~16'b0;
    assign data[5325] = ~16'b0;
    assign data[5326] = ~16'b0;
    assign data[5327] = ~16'b0;
    assign data[5328] = ~16'b0;
    assign data[5329] = ~16'b0;
    assign data[5330] = 16'b0;
    assign data[5331] = 16'b0;
    assign data[5332] = ~16'b0;
    assign data[5333] = ~16'b0;
    assign data[5334] = ~16'b0;
    assign data[5335] = ~16'b0;
    assign data[5336] = ~16'b0;
    assign data[5337] = ~16'b0;
    assign data[5338] = ~16'b0;
    assign data[5339] = ~16'b0;
    assign data[5340] = 16'b0;
    assign data[5341] = 16'b0;
    assign data[5342] = ~16'b0;
    assign data[5343] = ~16'b0;
    assign data[5344] = ~16'b0;
    assign data[5345] = ~16'b0;
    assign data[5346] = ~16'b0;
    assign data[5347] = ~16'b0;
    assign data[5348] = ~16'b0;
    assign data[5349] = ~16'b0;
    assign data[5350] = 16'b0;
    assign data[5351] = 16'b0;
    assign data[5352] = ~16'b0;
    assign data[5353] = ~16'b0;
    assign data[5354] = ~16'b0;
    assign data[5355] = ~16'b0;
    assign data[5356] = ~16'b0;
    assign data[5357] = ~16'b0;
    assign data[5358] = ~16'b0;
    assign data[5359] = ~16'b0;
    assign data[5360] = 16'b0;
    assign data[5361] = 16'b0;
    assign data[5362] = ~16'b0;
    assign data[5363] = ~16'b0;
    assign data[5364] = ~16'b0;
    assign data[5365] = ~16'b0;
    assign data[5366] = ~16'b0;
    assign data[5367] = ~16'b0;
    assign data[5368] = ~16'b0;
    assign data[5369] = ~16'b0;
    assign data[5370] = 16'b0;
    assign data[5371] = 16'b0;
    assign data[5372] = ~16'b0;
    assign data[5373] = ~16'b0;
    assign data[5374] = ~16'b0;
    assign data[5375] = ~16'b0;
    assign data[5376] = ~16'b0;
    assign data[5377] = ~16'b0;
    assign data[5378] = ~16'b0;
    assign data[5379] = ~16'b0;
    assign data[5380] = 16'b0;
    assign data[5381] = 16'b0;
    assign data[5382] = ~16'b0;
    assign data[5383] = ~16'b0;
    assign data[5384] = ~16'b0;
    assign data[5385] = ~16'b0;
    assign data[5386] = ~16'b0;
    assign data[5387] = ~16'b0;
    assign data[5388] = ~16'b0;
    assign data[5389] = ~16'b0;
    assign data[5390] = 16'b0;
    assign data[5391] = 16'b0;
    assign data[5392] = ~16'b0;
    assign data[5393] = ~16'b0;
    assign data[5394] = ~16'b0;
    assign data[5395] = ~16'b0;
    assign data[5396] = ~16'b0;
    assign data[5397] = ~16'b0;
    assign data[5398] = ~16'b0;
    assign data[5399] = ~16'b0;
    assign data[5400] = 16'b0;
    assign data[5401] = 16'b0;
    assign data[5402] = ~16'b0;
    assign data[5403] = ~16'b0;
    assign data[5404] = ~16'b0;
    assign data[5405] = ~16'b0;
    assign data[5406] = ~16'b0;
    assign data[5407] = ~16'b0;
    assign data[5408] = ~16'b0;
    assign data[5409] = ~16'b0;
    assign data[5410] = 16'b0;
    assign data[5411] = 16'b0;
    assign data[5412] = ~16'b0;
    assign data[5413] = ~16'b0;
    assign data[5414] = ~16'b0;
    assign data[5415] = ~16'b0;
    assign data[5416] = ~16'b0;
    assign data[5417] = ~16'b0;
    assign data[5418] = ~16'b0;
    assign data[5419] = ~16'b0;
    assign data[5420] = 16'b0;
    assign data[5421] = 16'b0;
    assign data[5422] = ~16'b0;
    assign data[5423] = ~16'b0;
    assign data[5424] = ~16'b0;
    assign data[5425] = ~16'b0;
    assign data[5426] = ~16'b0;
    assign data[5427] = ~16'b0;
    assign data[5428] = ~16'b0;
    assign data[5429] = ~16'b0;
    assign data[5430] = 16'b0;
    assign data[5431] = 16'b0;
    assign data[5432] = ~16'b0;
    assign data[5433] = ~16'b0;
    assign data[5434] = ~16'b0;
    assign data[5435] = ~16'b0;
    assign data[5436] = ~16'b0;
    assign data[5437] = ~16'b0;
    assign data[5438] = ~16'b0;
    assign data[5439] = ~16'b0;
    assign data[5440] = 16'b0;
    assign data[5441] = 16'b0;
    assign data[5442] = ~16'b0;
    assign data[5443] = ~16'b0;
    assign data[5444] = ~16'b0;
    assign data[5445] = ~16'b0;
    assign data[5446] = ~16'b0;
    assign data[5447] = ~16'b0;
    assign data[5448] = ~16'b0;
    assign data[5449] = ~16'b0;
    assign data[5450] = 16'b0;
    assign data[5451] = 16'b0;
    assign data[5452] = ~16'b0;
    assign data[5453] = ~16'b0;
    assign data[5454] = ~16'b0;
    assign data[5455] = ~16'b0;
    assign data[5456] = ~16'b0;
    assign data[5457] = ~16'b0;
    assign data[5458] = ~16'b0;
    assign data[5459] = ~16'b0;
    assign data[5460] = 16'b0;
    assign data[5461] = 16'b0;
    assign data[5462] = 16'b0;
    assign data[5463] = 16'b0;
    assign data[5464] = 16'b0;
    assign data[5465] = 16'b0;
    assign data[5466] = 16'b0;
    assign data[5467] = 16'b0;
    assign data[5468] = 16'b0;
    assign data[5469] = 16'b0;
    assign data[5470] = 16'b0;
    assign data[5471] = 16'b0;
    assign data[5472] = 16'b0;
    assign data[5473] = 16'b0;
    assign data[5474] = 16'b0;
    assign data[5475] = 16'b0;
    assign data[5476] = 16'b0;
    assign data[5477] = 16'b0;
    assign data[5478] = 16'b0;
    assign data[5479] = 16'b0;
    assign data[5480] = ~16'b0;
    assign data[5481] = ~16'b0;
    assign data[5482] = ~16'b0;
    assign data[5483] = ~16'b0;
    assign data[5484] = ~16'b0;
    assign data[5485] = ~16'b0;
    assign data[5486] = ~16'b0;
    assign data[5487] = ~16'b0;
    assign data[5488] = ~16'b0;
    assign data[5489] = ~16'b0;
    assign data[5490] = ~16'b0;
    assign data[5491] = ~16'b0;
    assign data[5492] = ~16'b0;
    assign data[5493] = ~16'b0;
    assign data[5494] = ~16'b0;
    assign data[5495] = ~16'b0;
    assign data[5496] = ~16'b0;
    assign data[5497] = ~16'b0;
    assign data[5498] = ~16'b0;
    assign data[5499] = ~16'b0;
    assign data[5500] = ~16'b0;
    assign data[5501] = ~16'b0;
    assign data[5502] = ~16'b0;
    assign data[5503] = ~16'b0;
    assign data[5504] = ~16'b0;
    assign data[5505] = ~16'b0;
    assign data[5506] = ~16'b0;
    assign data[5507] = ~16'b0;
    assign data[5508] = ~16'b0;
    assign data[5509] = ~16'b0;
    assign data[5510] = ~16'b0;
    assign data[5511] = ~16'b0;
    assign data[5512] = ~16'b0;
    assign data[5513] = ~16'b0;
    assign data[5514] = ~16'b0;
    assign data[5515] = ~16'b0;
    assign data[5516] = ~16'b0;
    assign data[5517] = ~16'b0;
    assign data[5518] = ~16'b0;
    assign data[5519] = ~16'b0;
    assign data[5520] = ~16'b0;
    assign data[5521] = ~16'b0;
    assign data[5522] = ~16'b0;
    assign data[5523] = ~16'b0;
    assign data[5524] = ~16'b0;
    assign data[5525] = ~16'b0;
    assign data[5526] = ~16'b0;
    assign data[5527] = ~16'b0;
    assign data[5528] = ~16'b0;
    assign data[5529] = ~16'b0;
    assign data[5530] = ~16'b0;
    assign data[5531] = ~16'b0;
    assign data[5532] = ~16'b0;
    assign data[5533] = ~16'b0;
    assign data[5534] = ~16'b0;
    assign data[5535] = ~16'b0;
    assign data[5536] = ~16'b0;
    assign data[5537] = ~16'b0;
    assign data[5538] = ~16'b0;
    assign data[5539] = ~16'b0;
    assign data[5540] = ~16'b0;
    assign data[5541] = ~16'b0;
    assign data[5542] = ~16'b0;
    assign data[5543] = ~16'b0;
    assign data[5544] = ~16'b0;
    assign data[5545] = ~16'b0;
    assign data[5546] = ~16'b0;
    assign data[5547] = ~16'b0;
    assign data[5548] = ~16'b0;
    assign data[5549] = ~16'b0;
    assign data[5550] = ~16'b0;
    assign data[5551] = ~16'b0;
    assign data[5552] = ~16'b0;
    assign data[5553] = ~16'b0;
    assign data[5554] = ~16'b0;
    assign data[5555] = ~16'b0;
    assign data[5556] = ~16'b0;
    assign data[5557] = ~16'b0;
    assign data[5558] = ~16'b0;
    assign data[5559] = ~16'b0;
    assign data[5560] = ~16'b0;
    assign data[5561] = ~16'b0;
    assign data[5562] = ~16'b0;
    assign data[5563] = ~16'b0;
    assign data[5564] = ~16'b0;
    assign data[5565] = ~16'b0;
    assign data[5566] = ~16'b0;
    assign data[5567] = ~16'b0;
    assign data[5568] = ~16'b0;
    assign data[5569] = ~16'b0;
    assign data[5570] = ~16'b0;
    assign data[5571] = ~16'b0;
    assign data[5572] = ~16'b0;
    assign data[5573] = ~16'b0;
    assign data[5574] = ~16'b0;
    assign data[5575] = ~16'b0;
    assign data[5576] = ~16'b0;
    assign data[5577] = ~16'b0;
    assign data[5578] = ~16'b0;
    assign data[5579] = ~16'b0;
    assign data[5580] = ~16'b0;
    assign data[5581] = ~16'b0;
    assign data[5582] = ~16'b0;
    assign data[5583] = ~16'b0;
    assign data[5584] = ~16'b0;
    assign data[5585] = ~16'b0;
    assign data[5586] = ~16'b0;
    assign data[5587] = ~16'b0;
    assign data[5588] = ~16'b0;
    assign data[5589] = ~16'b0;
    assign data[5590] = ~16'b0;
    assign data[5591] = ~16'b0;
    assign data[5592] = ~16'b0;
    assign data[5593] = ~16'b0;
    assign data[5594] = ~16'b0;
    assign data[5595] = ~16'b0;
    assign data[5596] = ~16'b0;
    assign data[5597] = ~16'b0;
    assign data[5598] = ~16'b0;
    assign data[5599] = ~16'b0;
    assign data[5600] = ~16'b0;
    assign data[5601] = ~16'b0;
    assign data[5602] = ~16'b0;
    assign data[5603] = ~16'b0;
    assign data[5604] = ~16'b0;
    assign data[5605] = ~16'b0;
    assign data[5606] = ~16'b0;
    assign data[5607] = ~16'b0;
    assign data[5608] = ~16'b0;
    assign data[5609] = ~16'b0;
    assign data[5610] = ~16'b0;
    assign data[5611] = ~16'b0;
    assign data[5612] = ~16'b0;
    assign data[5613] = ~16'b0;
    assign data[5614] = ~16'b0;
    assign data[5615] = ~16'b0;
    assign data[5616] = ~16'b0;
    assign data[5617] = ~16'b0;
    assign data[5618] = ~16'b0;
    assign data[5619] = ~16'b0;
    assign data[5620] = ~16'b0;
    assign data[5621] = ~16'b0;
    assign data[5622] = ~16'b0;
    assign data[5623] = ~16'b0;
    assign data[5624] = ~16'b0;
    assign data[5625] = ~16'b0;
    assign data[5626] = ~16'b0;
    assign data[5627] = ~16'b0;
    assign data[5628] = ~16'b0;
    assign data[5629] = ~16'b0;
    assign data[5630] = ~16'b0;
    assign data[5631] = ~16'b0;
    assign data[5632] = ~16'b0;
    assign data[5633] = ~16'b0;
    assign data[5634] = ~16'b0;
    assign data[5635] = ~16'b0;
    assign data[5636] = ~16'b0;
    assign data[5637] = ~16'b0;
    assign data[5638] = ~16'b0;
    assign data[5639] = ~16'b0;
    assign data[5640] = ~16'b0;
    assign data[5641] = ~16'b0;
    assign data[5642] = ~16'b0;
    assign data[5643] = ~16'b0;
    assign data[5644] = ~16'b0;
    assign data[5645] = ~16'b0;
    assign data[5646] = ~16'b0;
    assign data[5647] = ~16'b0;
    assign data[5648] = ~16'b0;
    assign data[5649] = ~16'b0;
    assign data[5650] = ~16'b0;
    assign data[5651] = ~16'b0;
    assign data[5652] = ~16'b0;
    assign data[5653] = ~16'b0;
    assign data[5654] = ~16'b0;
    assign data[5655] = ~16'b0;
    assign data[5656] = ~16'b0;
    assign data[5657] = ~16'b0;
    assign data[5658] = ~16'b0;
    assign data[5659] = ~16'b0;
    assign data[5660] = ~16'b0;
    assign data[5661] = ~16'b0;
    assign data[5662] = ~16'b0;
    assign data[5663] = ~16'b0;
    assign data[5664] = ~16'b0;
    assign data[5665] = ~16'b0;
    assign data[5666] = ~16'b0;
    assign data[5667] = ~16'b0;
    assign data[5668] = ~16'b0;
    assign data[5669] = ~16'b0;
    assign data[5670] = ~16'b0;
    assign data[5671] = ~16'b0;
    assign data[5672] = ~16'b0;
    assign data[5673] = ~16'b0;
    assign data[5674] = ~16'b0;
    assign data[5675] = ~16'b0;
    assign data[5676] = ~16'b0;
    assign data[5677] = ~16'b0;
    assign data[5678] = ~16'b0;
    assign data[5679] = ~16'b0;
    assign data[5680] = ~16'b0;
    assign data[5681] = ~16'b0;
    assign data[5682] = ~16'b0;
    assign data[5683] = ~16'b0;
    assign data[5684] = ~16'b0;
    assign data[5685] = ~16'b0;
    assign data[5686] = ~16'b0;
    assign data[5687] = ~16'b0;
    assign data[5688] = ~16'b0;
    assign data[5689] = ~16'b0;
    assign data[5690] = ~16'b0;
    assign data[5691] = ~16'b0;
    assign data[5692] = ~16'b0;
    assign data[5693] = ~16'b0;
    assign data[5694] = ~16'b0;
    assign data[5695] = ~16'b0;
    assign data[5696] = ~16'b0;
    assign data[5697] = ~16'b0;
    assign data[5698] = ~16'b0;
    assign data[5699] = ~16'b0;
    assign data[5700] = ~16'b0;
    assign data[5701] = ~16'b0;
    assign data[5702] = ~16'b0;
    assign data[5703] = ~16'b0;
    assign data[5704] = ~16'b0;
    assign data[5705] = ~16'b0;
    assign data[5706] = ~16'b0;
    assign data[5707] = ~16'b0;
    assign data[5708] = ~16'b0;
    assign data[5709] = ~16'b0;
    assign data[5710] = ~16'b0;
    assign data[5711] = ~16'b0;
    assign data[5712] = ~16'b0;
    assign data[5713] = ~16'b0;
    assign data[5714] = ~16'b0;
    assign data[5715] = ~16'b0;
    assign data[5716] = ~16'b0;
    assign data[5717] = ~16'b0;
    assign data[5718] = ~16'b0;
    assign data[5719] = ~16'b0;
    assign data[5720] = ~16'b0;
    assign data[5721] = ~16'b0;
    assign data[5722] = ~16'b0;
    assign data[5723] = ~16'b0;
    assign data[5724] = ~16'b0;
    assign data[5725] = ~16'b0;
    assign data[5726] = ~16'b0;
    assign data[5727] = ~16'b0;
    assign data[5728] = ~16'b0;
    assign data[5729] = ~16'b0;
    assign data[5730] = ~16'b0;
    assign data[5731] = ~16'b0;
    assign data[5732] = ~16'b0;
    assign data[5733] = ~16'b0;
    assign data[5734] = ~16'b0;
    assign data[5735] = ~16'b0;
    assign data[5736] = ~16'b0;
    assign data[5737] = ~16'b0;
    assign data[5738] = ~16'b0;
    assign data[5739] = ~16'b0;
    assign data[5740] = ~16'b0;
    assign data[5741] = ~16'b0;
    assign data[5742] = ~16'b0;
    assign data[5743] = ~16'b0;
    assign data[5744] = ~16'b0;
    assign data[5745] = ~16'b0;
    assign data[5746] = ~16'b0;
    assign data[5747] = ~16'b0;
    assign data[5748] = ~16'b0;
    assign data[5749] = ~16'b0;
    assign data[5750] = ~16'b0;
    assign data[5751] = ~16'b0;
    assign data[5752] = ~16'b0;
    assign data[5753] = ~16'b0;
    assign data[5754] = ~16'b0;
    assign data[5755] = ~16'b0;
    assign data[5756] = ~16'b0;
    assign data[5757] = ~16'b0;
    assign data[5758] = ~16'b0;
    assign data[5759] = ~16'b0;
    assign data[5760] = ~16'b0;
    assign data[5761] = ~16'b0;
    assign data[5762] = ~16'b0;
    assign data[5763] = ~16'b0;
    assign data[5764] = ~16'b0;
    assign data[5765] = ~16'b0;
    assign data[5766] = ~16'b0;
    assign data[5767] = ~16'b0;
    assign data[5768] = ~16'b0;
    assign data[5769] = ~16'b0;
    assign data[5770] = ~16'b0;
    assign data[5771] = ~16'b0;
    assign data[5772] = ~16'b0;
    assign data[5773] = ~16'b0;
    assign data[5774] = ~16'b0;
    assign data[5775] = ~16'b0;
    assign data[5776] = ~16'b0;
    assign data[5777] = ~16'b0;
    assign data[5778] = ~16'b0;
    assign data[5779] = ~16'b0;
    assign data[5780] = ~16'b0;
    assign data[5781] = ~16'b0;
    assign data[5782] = ~16'b0;
    assign data[5783] = ~16'b0;
    assign data[5784] = ~16'b0;
    assign data[5785] = ~16'b0;
    assign data[5786] = ~16'b0;
    assign data[5787] = ~16'b0;
    assign data[5788] = ~16'b0;
    assign data[5789] = ~16'b0;
    assign data[5790] = ~16'b0;
    assign data[5791] = ~16'b0;
    assign data[5792] = ~16'b0;
    assign data[5793] = ~16'b0;
    assign data[5794] = ~16'b0;
    assign data[5795] = ~16'b0;
    assign data[5796] = ~16'b0;
    assign data[5797] = ~16'b0;
    assign data[5798] = ~16'b0;
    assign data[5799] = ~16'b0;
    assign data[5800] = ~16'b0;
    assign data[5801] = ~16'b0;
    assign data[5802] = ~16'b0;
    assign data[5803] = ~16'b0;
    assign data[5804] = ~16'b0;
    assign data[5805] = ~16'b0;
    assign data[5806] = ~16'b0;
    assign data[5807] = ~16'b0;
    assign data[5808] = ~16'b0;
    assign data[5809] = ~16'b0;
    assign data[5810] = ~16'b0;
    assign data[5811] = ~16'b0;
    assign data[5812] = ~16'b0;
    assign data[5813] = ~16'b0;
    assign data[5814] = ~16'b0;
    assign data[5815] = ~16'b0;
    assign data[5816] = ~16'b0;
    assign data[5817] = ~16'b0;
    assign data[5818] = ~16'b0;
    assign data[5819] = ~16'b0;
    assign data[5820] = ~16'b0;
    assign data[5821] = ~16'b0;
    assign data[5822] = ~16'b0;
    assign data[5823] = ~16'b0;
    assign data[5824] = ~16'b0;
    assign data[5825] = ~16'b0;
    assign data[5826] = ~16'b0;
    assign data[5827] = ~16'b0;
    assign data[5828] = ~16'b0;
    assign data[5829] = ~16'b0;
    assign data[5830] = ~16'b0;
    assign data[5831] = ~16'b0;
    assign data[5832] = ~16'b0;
    assign data[5833] = ~16'b0;
    assign data[5834] = ~16'b0;
    assign data[5835] = ~16'b0;
    assign data[5836] = ~16'b0;
    assign data[5837] = ~16'b0;
    assign data[5838] = ~16'b0;
    assign data[5839] = ~16'b0;
    assign data[5840] = ~16'b0;
    assign data[5841] = ~16'b0;
    assign data[5842] = ~16'b0;
    assign data[5843] = ~16'b0;
    assign data[5844] = ~16'b0;
    assign data[5845] = ~16'b0;
    assign data[5846] = ~16'b0;
    assign data[5847] = ~16'b0;
    assign data[5848] = ~16'b0;
    assign data[5849] = ~16'b0;
    assign data[5850] = 16'b0;
    assign data[5851] = 16'b0;
    assign data[5852] = 16'b0;
    assign data[5853] = 16'b0;
    assign data[5854] = 16'b0;
    assign data[5855] = 16'b0;
    assign data[5856] = 16'b0;
    assign data[5857] = 16'b0;
    assign data[5858] = 16'b0;
    assign data[5859] = 16'b0;
    assign data[5860] = 16'b0;
    assign data[5861] = 16'b0;
    assign data[5862] = 16'b0;
    assign data[5863] = 16'b0;
    assign data[5864] = 16'b0;
    assign data[5865] = 16'b0;
    assign data[5866] = 16'b0;
    assign data[5867] = 16'b0;
    assign data[5868] = 16'b0;
    assign data[5869] = 16'b0;
    assign data[5870] = 16'b0;
    assign data[5871] = 16'b0;
    assign data[5872] = ~16'b0;
    assign data[5873] = ~16'b0;
    assign data[5874] = ~16'b0;
    assign data[5875] = ~16'b0;
    assign data[5876] = ~16'b0;
    assign data[5877] = ~16'b0;
    assign data[5878] = ~16'b0;
    assign data[5879] = ~16'b0;
    assign data[5880] = 16'b0;
    assign data[5881] = 16'b0;
    assign data[5882] = ~16'b0;
    assign data[5883] = ~16'b0;
    assign data[5884] = ~16'b0;
    assign data[5885] = ~16'b0;
    assign data[5886] = ~16'b0;
    assign data[5887] = ~16'b0;
    assign data[5888] = ~16'b0;
    assign data[5889] = ~16'b0;
    assign data[5890] = 16'b0;
    assign data[5891] = 16'b0;
    assign data[5892] = ~16'b0;
    assign data[5893] = ~16'b0;
    assign data[5894] = ~16'b0;
    assign data[5895] = ~16'b0;
    assign data[5896] = ~16'b0;
    assign data[5897] = ~16'b0;
    assign data[5898] = ~16'b0;
    assign data[5899] = ~16'b0;
    assign data[5900] = 16'b0;
    assign data[5901] = 16'b0;
    assign data[5902] = ~16'b0;
    assign data[5903] = ~16'b0;
    assign data[5904] = ~16'b0;
    assign data[5905] = ~16'b0;
    assign data[5906] = ~16'b0;
    assign data[5907] = ~16'b0;
    assign data[5908] = ~16'b0;
    assign data[5909] = ~16'b0;
    assign data[5910] = 16'b0;
    assign data[5911] = 16'b0;
    assign data[5912] = ~16'b0;
    assign data[5913] = ~16'b0;
    assign data[5914] = ~16'b0;
    assign data[5915] = ~16'b0;
    assign data[5916] = ~16'b0;
    assign data[5917] = ~16'b0;
    assign data[5918] = ~16'b0;
    assign data[5919] = ~16'b0;
    assign data[5920] = 16'b0;
    assign data[5921] = 16'b0;
    assign data[5922] = ~16'b0;
    assign data[5923] = ~16'b0;
    assign data[5924] = ~16'b0;
    assign data[5925] = ~16'b0;
    assign data[5926] = ~16'b0;
    assign data[5927] = ~16'b0;
    assign data[5928] = ~16'b0;
    assign data[5929] = ~16'b0;
    assign data[5930] = 16'b0;
    assign data[5931] = 16'b0;
    assign data[5932] = ~16'b0;
    assign data[5933] = ~16'b0;
    assign data[5934] = ~16'b0;
    assign data[5935] = ~16'b0;
    assign data[5936] = ~16'b0;
    assign data[5937] = ~16'b0;
    assign data[5938] = ~16'b0;
    assign data[5939] = ~16'b0;
    assign data[5940] = 16'b0;
    assign data[5941] = 16'b0;
    assign data[5942] = ~16'b0;
    assign data[5943] = ~16'b0;
    assign data[5944] = ~16'b0;
    assign data[5945] = ~16'b0;
    assign data[5946] = ~16'b0;
    assign data[5947] = ~16'b0;
    assign data[5948] = ~16'b0;
    assign data[5949] = ~16'b0;
    assign data[5950] = 16'b0;
    assign data[5951] = 16'b0;
    assign data[5952] = ~16'b0;
    assign data[5953] = ~16'b0;
    assign data[5954] = ~16'b0;
    assign data[5955] = ~16'b0;
    assign data[5956] = ~16'b0;
    assign data[5957] = ~16'b0;
    assign data[5958] = ~16'b0;
    assign data[5959] = ~16'b0;
    assign data[5960] = 16'b0;
    assign data[5961] = 16'b0;
    assign data[5962] = ~16'b0;
    assign data[5963] = ~16'b0;
    assign data[5964] = ~16'b0;
    assign data[5965] = ~16'b0;
    assign data[5966] = ~16'b0;
    assign data[5967] = ~16'b0;
    assign data[5968] = ~16'b0;
    assign data[5969] = ~16'b0;
    assign data[5970] = 16'b0;
    assign data[5971] = 16'b0;
    assign data[5972] = ~16'b0;
    assign data[5973] = ~16'b0;
    assign data[5974] = ~16'b0;
    assign data[5975] = ~16'b0;
    assign data[5976] = ~16'b0;
    assign data[5977] = ~16'b0;
    assign data[5978] = ~16'b0;
    assign data[5979] = ~16'b0;
    assign data[5980] = 16'b0;
    assign data[5981] = 16'b0;
    assign data[5982] = ~16'b0;
    assign data[5983] = ~16'b0;
    assign data[5984] = ~16'b0;
    assign data[5985] = ~16'b0;
    assign data[5986] = ~16'b0;
    assign data[5987] = ~16'b0;
    assign data[5988] = ~16'b0;
    assign data[5989] = ~16'b0;
    assign data[5990] = 16'b0;
    assign data[5991] = 16'b0;
    assign data[5992] = ~16'b0;
    assign data[5993] = ~16'b0;
    assign data[5994] = ~16'b0;
    assign data[5995] = ~16'b0;
    assign data[5996] = ~16'b0;
    assign data[5997] = ~16'b0;
    assign data[5998] = ~16'b0;
    assign data[5999] = ~16'b0;
    assign data[6000] = 16'b0;
    assign data[6001] = 16'b0;
    assign data[6002] = ~16'b0;
    assign data[6003] = ~16'b0;
    assign data[6004] = ~16'b0;
    assign data[6005] = ~16'b0;
    assign data[6006] = ~16'b0;
    assign data[6007] = ~16'b0;
    assign data[6008] = ~16'b0;
    assign data[6009] = ~16'b0;
    assign data[6010] = 16'b0;
    assign data[6011] = 16'b0;
    assign data[6012] = ~16'b0;
    assign data[6013] = ~16'b0;
    assign data[6014] = ~16'b0;
    assign data[6015] = ~16'b0;
    assign data[6016] = ~16'b0;
    assign data[6017] = ~16'b0;
    assign data[6018] = ~16'b0;
    assign data[6019] = ~16'b0;
    assign data[6020] = 16'b0;
    assign data[6021] = 16'b0;
    assign data[6022] = ~16'b0;
    assign data[6023] = ~16'b0;
    assign data[6024] = ~16'b0;
    assign data[6025] = ~16'b0;
    assign data[6026] = ~16'b0;
    assign data[6027] = ~16'b0;
    assign data[6028] = ~16'b0;
    assign data[6029] = ~16'b0;
    assign data[6030] = 16'b0;
    assign data[6031] = 16'b0;
    assign data[6032] = ~16'b0;
    assign data[6033] = ~16'b0;
    assign data[6034] = ~16'b0;
    assign data[6035] = ~16'b0;
    assign data[6036] = ~16'b0;
    assign data[6037] = ~16'b0;
    assign data[6038] = ~16'b0;
    assign data[6039] = ~16'b0;
    assign data[6040] = 16'b0;
    assign data[6041] = 16'b0;
    assign data[6042] = ~16'b0;
    assign data[6043] = ~16'b0;
    assign data[6044] = ~16'b0;
    assign data[6045] = ~16'b0;
    assign data[6046] = ~16'b0;
    assign data[6047] = ~16'b0;
    assign data[6048] = ~16'b0;
    assign data[6049] = ~16'b0;
    assign data[6050] = 16'b0;
    assign data[6051] = 16'b0;
    assign data[6052] = ~16'b0;
    assign data[6053] = ~16'b0;
    assign data[6054] = ~16'b0;
    assign data[6055] = ~16'b0;
    assign data[6056] = ~16'b0;
    assign data[6057] = ~16'b0;
    assign data[6058] = ~16'b0;
    assign data[6059] = ~16'b0;
    assign data[6060] = 16'b0;
    assign data[6061] = 16'b0;
    assign data[6062] = ~16'b0;
    assign data[6063] = ~16'b0;
    assign data[6064] = ~16'b0;
    assign data[6065] = ~16'b0;
    assign data[6066] = ~16'b0;
    assign data[6067] = ~16'b0;
    assign data[6068] = ~16'b0;
    assign data[6069] = ~16'b0;
    assign data[6070] = 16'b0;
    assign data[6071] = 16'b0;
    assign data[6072] = ~16'b0;
    assign data[6073] = ~16'b0;
    assign data[6074] = ~16'b0;
    assign data[6075] = ~16'b0;
    assign data[6076] = ~16'b0;
    assign data[6077] = ~16'b0;
    assign data[6078] = ~16'b0;
    assign data[6079] = ~16'b0;
    assign data[6080] = 16'b0;
    assign data[6081] = 16'b0;
    assign data[6082] = ~16'b0;
    assign data[6083] = ~16'b0;
    assign data[6084] = ~16'b0;
    assign data[6085] = ~16'b0;
    assign data[6086] = ~16'b0;
    assign data[6087] = ~16'b0;
    assign data[6088] = ~16'b0;
    assign data[6089] = ~16'b0;
    assign data[6090] = 16'b0;
    assign data[6091] = 16'b0;
    assign data[6092] = ~16'b0;
    assign data[6093] = ~16'b0;
    assign data[6094] = ~16'b0;
    assign data[6095] = ~16'b0;
    assign data[6096] = ~16'b0;
    assign data[6097] = ~16'b0;
    assign data[6098] = ~16'b0;
    assign data[6099] = ~16'b0;
    assign data[6100] = 16'b0;
    assign data[6101] = 16'b0;
    assign data[6102] = ~16'b0;
    assign data[6103] = ~16'b0;
    assign data[6104] = ~16'b0;
    assign data[6105] = ~16'b0;
    assign data[6106] = ~16'b0;
    assign data[6107] = ~16'b0;
    assign data[6108] = ~16'b0;
    assign data[6109] = ~16'b0;
    assign data[6110] = 16'b0;
    assign data[6111] = 16'b0;
    assign data[6112] = ~16'b0;
    assign data[6113] = ~16'b0;
    assign data[6114] = ~16'b0;
    assign data[6115] = ~16'b0;
    assign data[6116] = ~16'b0;
    assign data[6117] = ~16'b0;
    assign data[6118] = ~16'b0;
    assign data[6119] = ~16'b0;
    assign data[6120] = 16'b0;
    assign data[6121] = 16'b0;
    assign data[6122] = ~16'b0;
    assign data[6123] = ~16'b0;
    assign data[6124] = ~16'b0;
    assign data[6125] = ~16'b0;
    assign data[6126] = ~16'b0;
    assign data[6127] = ~16'b0;
    assign data[6128] = ~16'b0;
    assign data[6129] = ~16'b0;
    assign data[6130] = 16'b0;
    assign data[6131] = 16'b0;
    assign data[6132] = ~16'b0;
    assign data[6133] = ~16'b0;
    assign data[6134] = ~16'b0;
    assign data[6135] = ~16'b0;
    assign data[6136] = ~16'b0;
    assign data[6137] = ~16'b0;
    assign data[6138] = ~16'b0;
    assign data[6139] = ~16'b0;
    assign data[6140] = 16'b0;
    assign data[6141] = 16'b0;
    assign data[6142] = ~16'b0;
    assign data[6143] = ~16'b0;
    assign data[6144] = ~16'b0;
    assign data[6145] = ~16'b0;
    assign data[6146] = ~16'b0;
    assign data[6147] = ~16'b0;
    assign data[6148] = ~16'b0;
    assign data[6149] = ~16'b0;
    assign data[6150] = 16'b0;
    assign data[6151] = 16'b0;
    assign data[6152] = ~16'b0;
    assign data[6153] = ~16'b0;
    assign data[6154] = ~16'b0;
    assign data[6155] = ~16'b0;
    assign data[6156] = ~16'b0;
    assign data[6157] = ~16'b0;
    assign data[6158] = ~16'b0;
    assign data[6159] = ~16'b0;
    assign data[6160] = 16'b0;
    assign data[6161] = 16'b0;
    assign data[6162] = ~16'b0;
    assign data[6163] = ~16'b0;
    assign data[6164] = ~16'b0;
    assign data[6165] = ~16'b0;
    assign data[6166] = ~16'b0;
    assign data[6167] = ~16'b0;
    assign data[6168] = ~16'b0;
    assign data[6169] = ~16'b0;
    assign data[6170] = 16'b0;
    assign data[6171] = 16'b0;
    assign data[6172] = ~16'b0;
    assign data[6173] = ~16'b0;
    assign data[6174] = ~16'b0;
    assign data[6175] = ~16'b0;
    assign data[6176] = ~16'b0;
    assign data[6177] = ~16'b0;
    assign data[6178] = ~16'b0;
    assign data[6179] = ~16'b0;
    assign data[6180] = 16'b0;
    assign data[6181] = 16'b0;
    assign data[6182] = ~16'b0;
    assign data[6183] = ~16'b0;
    assign data[6184] = ~16'b0;
    assign data[6185] = ~16'b0;
    assign data[6186] = ~16'b0;
    assign data[6187] = ~16'b0;
    assign data[6188] = ~16'b0;
    assign data[6189] = ~16'b0;
    assign data[6190] = 16'b0;
    assign data[6191] = 16'b0;
    assign data[6192] = ~16'b0;
    assign data[6193] = ~16'b0;
    assign data[6194] = ~16'b0;
    assign data[6195] = ~16'b0;
    assign data[6196] = ~16'b0;
    assign data[6197] = ~16'b0;
    assign data[6198] = ~16'b0;
    assign data[6199] = ~16'b0;
    assign data[6200] = 16'b0;
    assign data[6201] = 16'b0;
    assign data[6202] = ~16'b0;
    assign data[6203] = ~16'b0;
    assign data[6204] = ~16'b0;
    assign data[6205] = ~16'b0;
    assign data[6206] = ~16'b0;
    assign data[6207] = ~16'b0;
    assign data[6208] = ~16'b0;
    assign data[6209] = ~16'b0;
    assign data[6210] = 16'b0;
    assign data[6211] = 16'b0;
    assign data[6212] = ~16'b0;
    assign data[6213] = ~16'b0;
    assign data[6214] = ~16'b0;
    assign data[6215] = ~16'b0;
    assign data[6216] = ~16'b0;
    assign data[6217] = ~16'b0;
    assign data[6218] = ~16'b0;
    assign data[6219] = ~16'b0;
    assign data[6220] = 16'b0;
    assign data[6221] = 16'b0;
    assign data[6222] = ~16'b0;
    assign data[6223] = ~16'b0;
    assign data[6224] = ~16'b0;
    assign data[6225] = ~16'b0;
    assign data[6226] = ~16'b0;
    assign data[6227] = ~16'b0;
    assign data[6228] = ~16'b0;
    assign data[6229] = ~16'b0;
    assign data[6230] = 16'b0;
    assign data[6231] = 16'b0;
    assign data[6232] = ~16'b0;
    assign data[6233] = ~16'b0;
    assign data[6234] = ~16'b0;
    assign data[6235] = ~16'b0;
    assign data[6236] = ~16'b0;
    assign data[6237] = ~16'b0;
    assign data[6238] = ~16'b0;
    assign data[6239] = ~16'b0;
    assign data[6240] = 16'b0;
    assign data[6241] = 16'b0;
    assign data[6242] = ~16'b0;
    assign data[6243] = ~16'b0;
    assign data[6244] = ~16'b0;
    assign data[6245] = ~16'b0;
    assign data[6246] = ~16'b0;
    assign data[6247] = ~16'b0;
    assign data[6248] = ~16'b0;
    assign data[6249] = ~16'b0;
    assign data[6250] = 16'b0;
    assign data[6251] = 16'b0;
    assign data[6252] = ~16'b0;
    assign data[6253] = ~16'b0;
    assign data[6254] = ~16'b0;
    assign data[6255] = ~16'b0;
    assign data[6256] = ~16'b0;
    assign data[6257] = ~16'b0;
    assign data[6258] = ~16'b0;
    assign data[6259] = ~16'b0;
    assign data[6260] = 16'b0;
    assign data[6261] = 16'b0;
    assign data[6262] = ~16'b0;
    assign data[6263] = ~16'b0;
    assign data[6264] = ~16'b0;
    assign data[6265] = ~16'b0;
    assign data[6266] = ~16'b0;
    assign data[6267] = ~16'b0;
    assign data[6268] = ~16'b0;
    assign data[6269] = ~16'b0;
    assign data[6270] = 16'b0;
    assign data[6271] = 16'b0;
    assign data[6272] = 16'b0;
    assign data[6273] = 16'b0;
    assign data[6274] = 16'b0;
    assign data[6275] = 16'b0;
    assign data[6276] = 16'b0;
    assign data[6277] = 16'b0;
    assign data[6278] = 16'b0;
    assign data[6279] = 16'b0;
    assign data[6280] = 16'b0;
    assign data[6281] = 16'b0;
    assign data[6282] = 16'b0;
    assign data[6283] = 16'b0;
    assign data[6284] = 16'b0;
    assign data[6285] = 16'b0;
    assign data[6286] = 16'b0;
    assign data[6287] = 16'b0;
    assign data[6288] = 16'b0;
    assign data[6289] = 16'b0;
    assign data[6290] = ~16'b0;
    assign data[6291] = ~16'b0;
    assign data[6292] = ~16'b0;
    assign data[6293] = ~16'b0;
    assign data[6294] = ~16'b0;
    assign data[6295] = ~16'b0;
    assign data[6296] = ~16'b0;
    assign data[6297] = ~16'b0;
    assign data[6298] = ~16'b0;
    assign data[6299] = ~16'b0;
    assign data[6300] = ~16'b0;
    assign data[6301] = ~16'b0;
    assign data[6302] = ~16'b0;
    assign data[6303] = ~16'b0;
    assign data[6304] = ~16'b0;
    assign data[6305] = ~16'b0;
    assign data[6306] = ~16'b0;
    assign data[6307] = ~16'b0;
    assign data[6308] = ~16'b0;
    assign data[6309] = ~16'b0;
    assign data[6310] = ~16'b0;
    assign data[6311] = ~16'b0;
    assign data[6312] = ~16'b0;
    assign data[6313] = ~16'b0;
    assign data[6314] = ~16'b0;
    assign data[6315] = ~16'b0;
    assign data[6316] = ~16'b0;
    assign data[6317] = ~16'b0;
    assign data[6318] = ~16'b0;
    assign data[6319] = ~16'b0;
    assign data[6320] = ~16'b0;
    assign data[6321] = ~16'b0;
    assign data[6322] = ~16'b0;
    assign data[6323] = ~16'b0;
    assign data[6324] = ~16'b0;
    assign data[6325] = ~16'b0;
    assign data[6326] = ~16'b0;
    assign data[6327] = ~16'b0;
    assign data[6328] = ~16'b0;
    assign data[6329] = ~16'b0;
    assign data[6330] = ~16'b0;
    assign data[6331] = ~16'b0;
    assign data[6332] = ~16'b0;
    assign data[6333] = ~16'b0;
    assign data[6334] = ~16'b0;
    assign data[6335] = ~16'b0;
    assign data[6336] = ~16'b0;
    assign data[6337] = ~16'b0;
    assign data[6338] = ~16'b0;
    assign data[6339] = ~16'b0;
    assign data[6340] = ~16'b0;
    assign data[6341] = ~16'b0;
    assign data[6342] = ~16'b0;
    assign data[6343] = ~16'b0;
    assign data[6344] = ~16'b0;
    assign data[6345] = ~16'b0;
    assign data[6346] = ~16'b0;
    assign data[6347] = ~16'b0;
    assign data[6348] = ~16'b0;
    assign data[6349] = ~16'b0;
    assign data[6350] = ~16'b0;
    assign data[6351] = ~16'b0;
    assign data[6352] = ~16'b0;
    assign data[6353] = ~16'b0;
    assign data[6354] = ~16'b0;
    assign data[6355] = ~16'b0;
    assign data[6356] = ~16'b0;
    assign data[6357] = ~16'b0;
    assign data[6358] = ~16'b0;
    assign data[6359] = ~16'b0;
    assign data[6360] = ~16'b0;
    assign data[6361] = ~16'b0;
    assign data[6362] = ~16'b0;
    assign data[6363] = ~16'b0;
    assign data[6364] = ~16'b0;
    assign data[6365] = ~16'b0;
    assign data[6366] = ~16'b0;
    assign data[6367] = ~16'b0;
    assign data[6368] = ~16'b0;
    assign data[6369] = ~16'b0;
    assign data[6370] = ~16'b0;
    assign data[6371] = ~16'b0;
    assign data[6372] = ~16'b0;
    assign data[6373] = ~16'b0;
    assign data[6374] = ~16'b0;
    assign data[6375] = ~16'b0;
    assign data[6376] = ~16'b0;
    assign data[6377] = ~16'b0;
    assign data[6378] = ~16'b0;
    assign data[6379] = ~16'b0;
    assign data[6380] = ~16'b0;
    assign data[6381] = ~16'b0;
    assign data[6382] = ~16'b0;
    assign data[6383] = ~16'b0;
    assign data[6384] = ~16'b0;
    assign data[6385] = ~16'b0;
    assign data[6386] = ~16'b0;
    assign data[6387] = ~16'b0;
    assign data[6388] = ~16'b0;
    assign data[6389] = ~16'b0;
    assign data[6390] = ~16'b0;
    assign data[6391] = ~16'b0;
    assign data[6392] = ~16'b0;
    assign data[6393] = ~16'b0;
    assign data[6394] = ~16'b0;
    assign data[6395] = ~16'b0;
    assign data[6396] = ~16'b0;
    assign data[6397] = ~16'b0;
    assign data[6398] = ~16'b0;
    assign data[6399] = ~16'b0;
    assign data[6400] = ~16'b0;
    assign data[6401] = ~16'b0;
    assign data[6402] = ~16'b0;
    assign data[6403] = ~16'b0;
    assign data[6404] = ~16'b0;
    assign data[6405] = ~16'b0;
    assign data[6406] = ~16'b0;
    assign data[6407] = ~16'b0;
    assign data[6408] = ~16'b0;
    assign data[6409] = ~16'b0;
    assign data[6410] = ~16'b0;
    assign data[6411] = ~16'b0;
    assign data[6412] = ~16'b0;
    assign data[6413] = ~16'b0;
    assign data[6414] = ~16'b0;
    assign data[6415] = ~16'b0;
    assign data[6416] = ~16'b0;
    assign data[6417] = ~16'b0;
    assign data[6418] = ~16'b0;
    assign data[6419] = ~16'b0;
    assign data[6420] = ~16'b0;
    assign data[6421] = ~16'b0;
    assign data[6422] = ~16'b0;
    assign data[6423] = ~16'b0;
    assign data[6424] = ~16'b0;
    assign data[6425] = ~16'b0;
    assign data[6426] = ~16'b0;
    assign data[6427] = ~16'b0;
    assign data[6428] = ~16'b0;
    assign data[6429] = ~16'b0;
    assign data[6430] = ~16'b0;
    assign data[6431] = ~16'b0;
    assign data[6432] = ~16'b0;
    assign data[6433] = ~16'b0;
    assign data[6434] = ~16'b0;
    assign data[6435] = ~16'b0;
    assign data[6436] = ~16'b0;
    assign data[6437] = ~16'b0;
    assign data[6438] = ~16'b0;
    assign data[6439] = ~16'b0;
    assign data[6440] = ~16'b0;
    assign data[6441] = ~16'b0;
    assign data[6442] = ~16'b0;
    assign data[6443] = ~16'b0;
    assign data[6444] = ~16'b0;
    assign data[6445] = ~16'b0;
    assign data[6446] = ~16'b0;
    assign data[6447] = ~16'b0;
    assign data[6448] = ~16'b0;
    assign data[6449] = ~16'b0;
    assign data[6450] = ~16'b0;
    assign data[6451] = ~16'b0;
    assign data[6452] = ~16'b0;
    assign data[6453] = ~16'b0;
    assign data[6454] = ~16'b0;
    assign data[6455] = ~16'b0;
    assign data[6456] = ~16'b0;
    assign data[6457] = ~16'b0;
    assign data[6458] = ~16'b0;
    assign data[6459] = ~16'b0;
    assign data[6460] = ~16'b0;
    assign data[6461] = ~16'b0;
    assign data[6462] = ~16'b0;
    assign data[6463] = ~16'b0;
    assign data[6464] = ~16'b0;
    assign data[6465] = ~16'b0;
    assign data[6466] = ~16'b0;
    assign data[6467] = ~16'b0;
    assign data[6468] = ~16'b0;
    assign data[6469] = ~16'b0;
    assign data[6470] = ~16'b0;
    assign data[6471] = ~16'b0;
    assign data[6472] = ~16'b0;
    assign data[6473] = ~16'b0;
    assign data[6474] = ~16'b0;
    assign data[6475] = ~16'b0;
    assign data[6476] = ~16'b0;
    assign data[6477] = ~16'b0;
    assign data[6478] = ~16'b0;
    assign data[6479] = ~16'b0;
    assign data[6480] = ~16'b0;
    assign data[6481] = ~16'b0;
    assign data[6482] = ~16'b0;
    assign data[6483] = ~16'b0;
    assign data[6484] = ~16'b0;
    assign data[6485] = ~16'b0;
    assign data[6486] = ~16'b0;
    assign data[6487] = ~16'b0;
    assign data[6488] = ~16'b0;
    assign data[6489] = ~16'b0;
    assign data[6490] = ~16'b0;
    assign data[6491] = ~16'b0;
    assign data[6492] = ~16'b0;
    assign data[6493] = ~16'b0;
    assign data[6494] = ~16'b0;
    assign data[6495] = ~16'b0;
    assign data[6496] = ~16'b0;
    assign data[6497] = ~16'b0;
    assign data[6498] = ~16'b0;
    assign data[6499] = ~16'b0;
    assign data[6500] = ~16'b0;
    assign data[6501] = ~16'b0;
    assign data[6502] = ~16'b0;
    assign data[6503] = ~16'b0;
    assign data[6504] = ~16'b0;
    assign data[6505] = ~16'b0;
    assign data[6506] = ~16'b0;
    assign data[6507] = ~16'b0;
    assign data[6508] = ~16'b0;
    assign data[6509] = ~16'b0;
    assign data[6510] = ~16'b0;
    assign data[6511] = ~16'b0;
    assign data[6512] = ~16'b0;
    assign data[6513] = ~16'b0;
    assign data[6514] = ~16'b0;
    assign data[6515] = ~16'b0;
    assign data[6516] = ~16'b0;
    assign data[6517] = ~16'b0;
    assign data[6518] = ~16'b0;
    assign data[6519] = ~16'b0;
    assign data[6520] = ~16'b0;
    assign data[6521] = ~16'b0;
    assign data[6522] = ~16'b0;
    assign data[6523] = ~16'b0;
    assign data[6524] = ~16'b0;
    assign data[6525] = ~16'b0;
    assign data[6526] = ~16'b0;
    assign data[6527] = ~16'b0;
    assign data[6528] = ~16'b0;
    assign data[6529] = ~16'b0;
    assign data[6530] = ~16'b0;
    assign data[6531] = ~16'b0;
    assign data[6532] = ~16'b0;
    assign data[6533] = ~16'b0;
    assign data[6534] = ~16'b0;
    assign data[6535] = ~16'b0;
    assign data[6536] = ~16'b0;
    assign data[6537] = ~16'b0;
    assign data[6538] = ~16'b0;
    assign data[6539] = ~16'b0;
    assign data[6540] = ~16'b0;
    assign data[6541] = ~16'b0;
    assign data[6542] = ~16'b0;
    assign data[6543] = ~16'b0;
    assign data[6544] = ~16'b0;
    assign data[6545] = ~16'b0;
    assign data[6546] = ~16'b0;
    assign data[6547] = ~16'b0;
    assign data[6548] = ~16'b0;
    assign data[6549] = ~16'b0;
    assign data[6550] = ~16'b0;
    assign data[6551] = ~16'b0;
    assign data[6552] = ~16'b0;
    assign data[6553] = ~16'b0;
    assign data[6554] = ~16'b0;
    assign data[6555] = ~16'b0;
    assign data[6556] = ~16'b0;
    assign data[6557] = ~16'b0;
    assign data[6558] = ~16'b0;
    assign data[6559] = ~16'b0;
    assign data[6560] = ~16'b0;
    assign data[6561] = ~16'b0;
    assign data[6562] = ~16'b0;
    assign data[6563] = ~16'b0;
    assign data[6564] = ~16'b0;
    assign data[6565] = ~16'b0;
    assign data[6566] = ~16'b0;
    assign data[6567] = ~16'b0;
    assign data[6568] = ~16'b0;
    assign data[6569] = ~16'b0;
    assign data[6570] = ~16'b0;
    assign data[6571] = ~16'b0;
    assign data[6572] = ~16'b0;
    assign data[6573] = ~16'b0;
    assign data[6574] = ~16'b0;
    assign data[6575] = ~16'b0;
    assign data[6576] = ~16'b0;
    assign data[6577] = ~16'b0;
    assign data[6578] = ~16'b0;
    assign data[6579] = ~16'b0;
    assign data[6580] = ~16'b0;
    assign data[6581] = ~16'b0;
    assign data[6582] = ~16'b0;
    assign data[6583] = ~16'b0;
    assign data[6584] = ~16'b0;
    assign data[6585] = ~16'b0;
    assign data[6586] = ~16'b0;
    assign data[6587] = ~16'b0;
    assign data[6588] = ~16'b0;
    assign data[6589] = ~16'b0;
    assign data[6590] = ~16'b0;
    assign data[6591] = ~16'b0;
    assign data[6592] = ~16'b0;
    assign data[6593] = ~16'b0;
    assign data[6594] = ~16'b0;
    assign data[6595] = ~16'b0;
    assign data[6596] = ~16'b0;
    assign data[6597] = ~16'b0;
    assign data[6598] = ~16'b0;
    assign data[6599] = ~16'b0;
    assign data[6600] = ~16'b0;
    assign data[6601] = ~16'b0;
    assign data[6602] = ~16'b0;
    assign data[6603] = ~16'b0;
    assign data[6604] = ~16'b0;
    assign data[6605] = ~16'b0;
    assign data[6606] = ~16'b0;
    assign data[6607] = ~16'b0;
    assign data[6608] = ~16'b0;
    assign data[6609] = ~16'b0;
    assign data[6610] = ~16'b0;
    assign data[6611] = ~16'b0;
    assign data[6612] = ~16'b0;
    assign data[6613] = ~16'b0;
    assign data[6614] = ~16'b0;
    assign data[6615] = ~16'b0;
    assign data[6616] = ~16'b0;
    assign data[6617] = ~16'b0;
    assign data[6618] = ~16'b0;
    assign data[6619] = ~16'b0;
    assign data[6620] = ~16'b0;
    assign data[6621] = ~16'b0;
    assign data[6622] = ~16'b0;
    assign data[6623] = ~16'b0;
    assign data[6624] = ~16'b0;
    assign data[6625] = ~16'b0;
    assign data[6626] = ~16'b0;
    assign data[6627] = ~16'b0;
    assign data[6628] = ~16'b0;
    assign data[6629] = ~16'b0;
    assign data[6630] = ~16'b0;
    assign data[6631] = ~16'b0;
    assign data[6632] = ~16'b0;
    assign data[6633] = ~16'b0;
    assign data[6634] = ~16'b0;
    assign data[6635] = ~16'b0;
    assign data[6636] = ~16'b0;
    assign data[6637] = ~16'b0;
    assign data[6638] = ~16'b0;
    assign data[6639] = ~16'b0;
    assign data[6640] = ~16'b0;
    assign data[6641] = ~16'b0;
    assign data[6642] = ~16'b0;
    assign data[6643] = ~16'b0;
    assign data[6644] = ~16'b0;
    assign data[6645] = ~16'b0;
    assign data[6646] = ~16'b0;
    assign data[6647] = ~16'b0;
    assign data[6648] = ~16'b0;
    assign data[6649] = ~16'b0;
    assign data[6650] = ~16'b0;
    assign data[6651] = ~16'b0;
    assign data[6652] = ~16'b0;
    assign data[6653] = ~16'b0;
    assign data[6654] = ~16'b0;
    assign data[6655] = ~16'b0;
    assign data[6656] = ~16'b0;
    assign data[6657] = ~16'b0;
    assign data[6658] = ~16'b0;
    assign data[6659] = ~16'b0;
    assign data[6660] = 16'b0;
    assign data[6661] = 16'b0;
    assign data[6662] = 16'b0;
    assign data[6663] = 16'b0;
    assign data[6664] = 16'b0;
    assign data[6665] = 16'b0;
    assign data[6666] = 16'b0;
    assign data[6667] = 16'b0;
    assign data[6668] = 16'b0;
    assign data[6669] = 16'b0;
    assign data[6670] = 16'b0;
    assign data[6671] = 16'b0;
    assign data[6672] = 16'b0;
    assign data[6673] = 16'b0;
    assign data[6674] = 16'b0;
    assign data[6675] = 16'b0;
    assign data[6676] = 16'b0;
    assign data[6677] = 16'b0;
    assign data[6678] = 16'b0;
    assign data[6679] = 16'b0;
    assign data[6680] = 16'b0;
    assign data[6681] = 16'b0;
    assign data[6682] = ~16'b0;
    assign data[6683] = ~16'b0;
    assign data[6684] = ~16'b0;
    assign data[6685] = ~16'b0;
    assign data[6686] = ~16'b0;
    assign data[6687] = ~16'b0;
    assign data[6688] = ~16'b0;
    assign data[6689] = ~16'b0;
    assign data[6690] = 16'b0;
    assign data[6691] = 16'b0;
    assign data[6692] = ~16'b0;
    assign data[6693] = ~16'b0;
    assign data[6694] = ~16'b0;
    assign data[6695] = ~16'b0;
    assign data[6696] = ~16'b0;
    assign data[6697] = ~16'b0;
    assign data[6698] = ~16'b0;
    assign data[6699] = ~16'b0;
    assign data[6700] = 16'b0;
    assign data[6701] = 16'b0;
    assign data[6702] = ~16'b0;
    assign data[6703] = ~16'b0;
    assign data[6704] = ~16'b0;
    assign data[6705] = ~16'b0;
    assign data[6706] = ~16'b0;
    assign data[6707] = ~16'b0;
    assign data[6708] = ~16'b0;
    assign data[6709] = ~16'b0;
    assign data[6710] = 16'b0;
    assign data[6711] = 16'b0;
    assign data[6712] = ~16'b0;
    assign data[6713] = ~16'b0;
    assign data[6714] = ~16'b0;
    assign data[6715] = ~16'b0;
    assign data[6716] = ~16'b0;
    assign data[6717] = ~16'b0;
    assign data[6718] = ~16'b0;
    assign data[6719] = ~16'b0;
    assign data[6720] = 16'b0;
    assign data[6721] = 16'b0;
    assign data[6722] = ~16'b0;
    assign data[6723] = ~16'b0;
    assign data[6724] = ~16'b0;
    assign data[6725] = ~16'b0;
    assign data[6726] = ~16'b0;
    assign data[6727] = ~16'b0;
    assign data[6728] = ~16'b0;
    assign data[6729] = ~16'b0;
    assign data[6730] = 16'b0;
    assign data[6731] = 16'b0;
    assign data[6732] = ~16'b0;
    assign data[6733] = ~16'b0;
    assign data[6734] = ~16'b0;
    assign data[6735] = ~16'b0;
    assign data[6736] = ~16'b0;
    assign data[6737] = ~16'b0;
    assign data[6738] = ~16'b0;
    assign data[6739] = ~16'b0;
    assign data[6740] = 16'b0;
    assign data[6741] = 16'b0;
    assign data[6742] = ~16'b0;
    assign data[6743] = ~16'b0;
    assign data[6744] = ~16'b0;
    assign data[6745] = ~16'b0;
    assign data[6746] = ~16'b0;
    assign data[6747] = ~16'b0;
    assign data[6748] = ~16'b0;
    assign data[6749] = ~16'b0;
    assign data[6750] = 16'b0;
    assign data[6751] = 16'b0;
    assign data[6752] = ~16'b0;
    assign data[6753] = ~16'b0;
    assign data[6754] = ~16'b0;
    assign data[6755] = ~16'b0;
    assign data[6756] = ~16'b0;
    assign data[6757] = ~16'b0;
    assign data[6758] = ~16'b0;
    assign data[6759] = ~16'b0;
    assign data[6760] = 16'b0;
    assign data[6761] = 16'b0;
    assign data[6762] = ~16'b0;
    assign data[6763] = ~16'b0;
    assign data[6764] = ~16'b0;
    assign data[6765] = ~16'b0;
    assign data[6766] = ~16'b0;
    assign data[6767] = ~16'b0;
    assign data[6768] = ~16'b0;
    assign data[6769] = ~16'b0;
    assign data[6770] = 16'b0;
    assign data[6771] = 16'b0;
    assign data[6772] = ~16'b0;
    assign data[6773] = ~16'b0;
    assign data[6774] = ~16'b0;
    assign data[6775] = ~16'b0;
    assign data[6776] = ~16'b0;
    assign data[6777] = ~16'b0;
    assign data[6778] = ~16'b0;
    assign data[6779] = ~16'b0;
    assign data[6780] = 16'b0;
    assign data[6781] = 16'b0;
    assign data[6782] = ~16'b0;
    assign data[6783] = ~16'b0;
    assign data[6784] = ~16'b0;
    assign data[6785] = ~16'b0;
    assign data[6786] = ~16'b0;
    assign data[6787] = ~16'b0;
    assign data[6788] = ~16'b0;
    assign data[6789] = ~16'b0;
    assign data[6790] = 16'b0;
    assign data[6791] = 16'b0;
    assign data[6792] = ~16'b0;
    assign data[6793] = ~16'b0;
    assign data[6794] = ~16'b0;
    assign data[6795] = ~16'b0;
    assign data[6796] = ~16'b0;
    assign data[6797] = ~16'b0;
    assign data[6798] = ~16'b0;
    assign data[6799] = ~16'b0;
    assign data[6800] = 16'b0;
    assign data[6801] = 16'b0;
    assign data[6802] = ~16'b0;
    assign data[6803] = ~16'b0;
    assign data[6804] = ~16'b0;
    assign data[6805] = ~16'b0;
    assign data[6806] = ~16'b0;
    assign data[6807] = ~16'b0;
    assign data[6808] = ~16'b0;
    assign data[6809] = ~16'b0;
    assign data[6810] = 16'b0;
    assign data[6811] = 16'b0;
    assign data[6812] = ~16'b0;
    assign data[6813] = ~16'b0;
    assign data[6814] = ~16'b0;
    assign data[6815] = ~16'b0;
    assign data[6816] = ~16'b0;
    assign data[6817] = ~16'b0;
    assign data[6818] = ~16'b0;
    assign data[6819] = ~16'b0;
    assign data[6820] = 16'b0;
    assign data[6821] = 16'b0;
    assign data[6822] = ~16'b0;
    assign data[6823] = ~16'b0;
    assign data[6824] = ~16'b0;
    assign data[6825] = ~16'b0;
    assign data[6826] = ~16'b0;
    assign data[6827] = ~16'b0;
    assign data[6828] = ~16'b0;
    assign data[6829] = ~16'b0;
    assign data[6830] = 16'b0;
    assign data[6831] = 16'b0;
    assign data[6832] = ~16'b0;
    assign data[6833] = ~16'b0;
    assign data[6834] = ~16'b0;
    assign data[6835] = ~16'b0;
    assign data[6836] = ~16'b0;
    assign data[6837] = ~16'b0;
    assign data[6838] = ~16'b0;
    assign data[6839] = ~16'b0;
    assign data[6840] = 16'b0;
    assign data[6841] = 16'b0;
    assign data[6842] = ~16'b0;
    assign data[6843] = ~16'b0;
    assign data[6844] = ~16'b0;
    assign data[6845] = ~16'b0;
    assign data[6846] = ~16'b0;
    assign data[6847] = ~16'b0;
    assign data[6848] = ~16'b0;
    assign data[6849] = ~16'b0;
    assign data[6850] = 16'b0;
    assign data[6851] = 16'b0;
    assign data[6852] = ~16'b0;
    assign data[6853] = ~16'b0;
    assign data[6854] = ~16'b0;
    assign data[6855] = ~16'b0;
    assign data[6856] = ~16'b0;
    assign data[6857] = ~16'b0;
    assign data[6858] = ~16'b0;
    assign data[6859] = ~16'b0;
    assign data[6860] = 16'b0;
    assign data[6861] = 16'b0;
    assign data[6862] = ~16'b0;
    assign data[6863] = ~16'b0;
    assign data[6864] = ~16'b0;
    assign data[6865] = ~16'b0;
    assign data[6866] = ~16'b0;
    assign data[6867] = ~16'b0;
    assign data[6868] = ~16'b0;
    assign data[6869] = ~16'b0;
    assign data[6870] = 16'b0;
    assign data[6871] = 16'b0;
    assign data[6872] = ~16'b0;
    assign data[6873] = ~16'b0;
    assign data[6874] = ~16'b0;
    assign data[6875] = ~16'b0;
    assign data[6876] = ~16'b0;
    assign data[6877] = ~16'b0;
    assign data[6878] = ~16'b0;
    assign data[6879] = ~16'b0;
    assign data[6880] = 16'b0;
    assign data[6881] = 16'b0;
    assign data[6882] = ~16'b0;
    assign data[6883] = ~16'b0;
    assign data[6884] = ~16'b0;
    assign data[6885] = ~16'b0;
    assign data[6886] = ~16'b0;
    assign data[6887] = ~16'b0;
    assign data[6888] = ~16'b0;
    assign data[6889] = ~16'b0;
    assign data[6890] = 16'b0;
    assign data[6891] = 16'b0;
    assign data[6892] = ~16'b0;
    assign data[6893] = ~16'b0;
    assign data[6894] = ~16'b0;
    assign data[6895] = ~16'b0;
    assign data[6896] = ~16'b0;
    assign data[6897] = ~16'b0;
    assign data[6898] = ~16'b0;
    assign data[6899] = ~16'b0;
    assign data[6900] = 16'b0;
    assign data[6901] = 16'b0;
    assign data[6902] = ~16'b0;
    assign data[6903] = ~16'b0;
    assign data[6904] = ~16'b0;
    assign data[6905] = ~16'b0;
    assign data[6906] = ~16'b0;
    assign data[6907] = ~16'b0;
    assign data[6908] = ~16'b0;
    assign data[6909] = ~16'b0;
    assign data[6910] = 16'b0;
    assign data[6911] = 16'b0;
    assign data[6912] = ~16'b0;
    assign data[6913] = ~16'b0;
    assign data[6914] = ~16'b0;
    assign data[6915] = ~16'b0;
    assign data[6916] = ~16'b0;
    assign data[6917] = ~16'b0;
    assign data[6918] = ~16'b0;
    assign data[6919] = ~16'b0;
    assign data[6920] = 16'b0;
    assign data[6921] = 16'b0;
    assign data[6922] = ~16'b0;
    assign data[6923] = ~16'b0;
    assign data[6924] = ~16'b0;
    assign data[6925] = ~16'b0;
    assign data[6926] = ~16'b0;
    assign data[6927] = ~16'b0;
    assign data[6928] = ~16'b0;
    assign data[6929] = ~16'b0;
    assign data[6930] = 16'b0;
    assign data[6931] = 16'b0;
    assign data[6932] = ~16'b0;
    assign data[6933] = ~16'b0;
    assign data[6934] = ~16'b0;
    assign data[6935] = ~16'b0;
    assign data[6936] = ~16'b0;
    assign data[6937] = ~16'b0;
    assign data[6938] = ~16'b0;
    assign data[6939] = ~16'b0;
    assign data[6940] = 16'b0;
    assign data[6941] = 16'b0;
    assign data[6942] = ~16'b0;
    assign data[6943] = ~16'b0;
    assign data[6944] = ~16'b0;
    assign data[6945] = ~16'b0;
    assign data[6946] = ~16'b0;
    assign data[6947] = ~16'b0;
    assign data[6948] = ~16'b0;
    assign data[6949] = ~16'b0;
    assign data[6950] = 16'b0;
    assign data[6951] = 16'b0;
    assign data[6952] = ~16'b0;
    assign data[6953] = ~16'b0;
    assign data[6954] = ~16'b0;
    assign data[6955] = ~16'b0;
    assign data[6956] = ~16'b0;
    assign data[6957] = ~16'b0;
    assign data[6958] = ~16'b0;
    assign data[6959] = ~16'b0;
    assign data[6960] = 16'b0;
    assign data[6961] = 16'b0;
    assign data[6962] = ~16'b0;
    assign data[6963] = ~16'b0;
    assign data[6964] = ~16'b0;
    assign data[6965] = ~16'b0;
    assign data[6966] = ~16'b0;
    assign data[6967] = ~16'b0;
    assign data[6968] = ~16'b0;
    assign data[6969] = ~16'b0;
    assign data[6970] = 16'b0;
    assign data[6971] = 16'b0;
    assign data[6972] = ~16'b0;
    assign data[6973] = ~16'b0;
    assign data[6974] = ~16'b0;
    assign data[6975] = ~16'b0;
    assign data[6976] = ~16'b0;
    assign data[6977] = ~16'b0;
    assign data[6978] = ~16'b0;
    assign data[6979] = ~16'b0;
    assign data[6980] = 16'b0;
    assign data[6981] = 16'b0;
    assign data[6982] = ~16'b0;
    assign data[6983] = ~16'b0;
    assign data[6984] = ~16'b0;
    assign data[6985] = ~16'b0;
    assign data[6986] = ~16'b0;
    assign data[6987] = ~16'b0;
    assign data[6988] = ~16'b0;
    assign data[6989] = ~16'b0;
    assign data[6990] = 16'b0;
    assign data[6991] = 16'b0;
    assign data[6992] = ~16'b0;
    assign data[6993] = ~16'b0;
    assign data[6994] = ~16'b0;
    assign data[6995] = ~16'b0;
    assign data[6996] = ~16'b0;
    assign data[6997] = ~16'b0;
    assign data[6998] = ~16'b0;
    assign data[6999] = ~16'b0;
    assign data[7000] = 16'b0;
    assign data[7001] = 16'b0;
    assign data[7002] = ~16'b0;
    assign data[7003] = ~16'b0;
    assign data[7004] = ~16'b0;
    assign data[7005] = ~16'b0;
    assign data[7006] = ~16'b0;
    assign data[7007] = ~16'b0;
    assign data[7008] = ~16'b0;
    assign data[7009] = ~16'b0;
    assign data[7010] = 16'b0;
    assign data[7011] = 16'b0;
    assign data[7012] = ~16'b0;
    assign data[7013] = ~16'b0;
    assign data[7014] = ~16'b0;
    assign data[7015] = ~16'b0;
    assign data[7016] = ~16'b0;
    assign data[7017] = ~16'b0;
    assign data[7018] = ~16'b0;
    assign data[7019] = ~16'b0;
    assign data[7020] = 16'b0;
    assign data[7021] = 16'b0;
    assign data[7022] = ~16'b0;
    assign data[7023] = ~16'b0;
    assign data[7024] = ~16'b0;
    assign data[7025] = ~16'b0;
    assign data[7026] = ~16'b0;
    assign data[7027] = ~16'b0;
    assign data[7028] = ~16'b0;
    assign data[7029] = ~16'b0;
    assign data[7030] = 16'b0;
    assign data[7031] = 16'b0;
    assign data[7032] = ~16'b0;
    assign data[7033] = ~16'b0;
    assign data[7034] = ~16'b0;
    assign data[7035] = ~16'b0;
    assign data[7036] = ~16'b0;
    assign data[7037] = ~16'b0;
    assign data[7038] = ~16'b0;
    assign data[7039] = ~16'b0;
    assign data[7040] = 16'b0;
    assign data[7041] = 16'b0;
    assign data[7042] = ~16'b0;
    assign data[7043] = ~16'b0;
    assign data[7044] = ~16'b0;
    assign data[7045] = ~16'b0;
    assign data[7046] = ~16'b0;
    assign data[7047] = ~16'b0;
    assign data[7048] = ~16'b0;
    assign data[7049] = ~16'b0;
    assign data[7050] = 16'b0;
    assign data[7051] = 16'b0;
    assign data[7052] = ~16'b0;
    assign data[7053] = ~16'b0;
    assign data[7054] = ~16'b0;
    assign data[7055] = ~16'b0;
    assign data[7056] = ~16'b0;
    assign data[7057] = ~16'b0;
    assign data[7058] = ~16'b0;
    assign data[7059] = ~16'b0;
    assign data[7060] = 16'b0;
    assign data[7061] = 16'b0;
    assign data[7062] = ~16'b0;
    assign data[7063] = ~16'b0;
    assign data[7064] = ~16'b0;
    assign data[7065] = ~16'b0;
    assign data[7066] = ~16'b0;
    assign data[7067] = ~16'b0;
    assign data[7068] = ~16'b0;
    assign data[7069] = ~16'b0;
    assign data[7070] = 16'b0;
    assign data[7071] = 16'b0;
    assign data[7072] = ~16'b0;
    assign data[7073] = ~16'b0;
    assign data[7074] = ~16'b0;
    assign data[7075] = ~16'b0;
    assign data[7076] = ~16'b0;
    assign data[7077] = ~16'b0;
    assign data[7078] = ~16'b0;
    assign data[7079] = ~16'b0;
    assign data[7080] = 16'b0;
    assign data[7081] = 16'b0;
    assign data[7082] = 16'b0;
    assign data[7083] = 16'b0;
    assign data[7084] = 16'b0;
    assign data[7085] = 16'b0;
    assign data[7086] = 16'b0;
    assign data[7087] = 16'b0;
    assign data[7088] = 16'b0;
    assign data[7089] = 16'b0;
    assign data[7090] = 16'b0;
    assign data[7091] = 16'b0;
    assign data[7092] = 16'b0;
    assign data[7093] = 16'b0;
    assign data[7094] = 16'b0;
    assign data[7095] = 16'b0;
    assign data[7096] = 16'b0;
    assign data[7097] = 16'b0;
    assign data[7098] = 16'b0;
    assign data[7099] = 16'b0;
    assign data[7100] = ~16'b0;
    assign data[7101] = ~16'b0;
    assign data[7102] = ~16'b0;
    assign data[7103] = ~16'b0;
    assign data[7104] = ~16'b0;
    assign data[7105] = ~16'b0;
    assign data[7106] = ~16'b0;
    assign data[7107] = ~16'b0;
    assign data[7108] = ~16'b0;
    assign data[7109] = ~16'b0;
    assign data[7110] = ~16'b0;
    assign data[7111] = ~16'b0;
    assign data[7112] = ~16'b0;
    assign data[7113] = ~16'b0;
    assign data[7114] = ~16'b0;
    assign data[7115] = ~16'b0;
    assign data[7116] = ~16'b0;
    assign data[7117] = ~16'b0;
    assign data[7118] = ~16'b0;
    assign data[7119] = ~16'b0;
    assign data[7120] = ~16'b0;
    assign data[7121] = ~16'b0;
    assign data[7122] = ~16'b0;
    assign data[7123] = ~16'b0;
    assign data[7124] = ~16'b0;
    assign data[7125] = ~16'b0;
    assign data[7126] = ~16'b0;
    assign data[7127] = ~16'b0;
    assign data[7128] = ~16'b0;
    assign data[7129] = ~16'b0;
    assign data[7130] = ~16'b0;
    assign data[7131] = ~16'b0;
    assign data[7132] = ~16'b0;
    assign data[7133] = ~16'b0;
    assign data[7134] = ~16'b0;
    assign data[7135] = ~16'b0;
    assign data[7136] = ~16'b0;
    assign data[7137] = ~16'b0;
    assign data[7138] = ~16'b0;
    assign data[7139] = ~16'b0;
    assign data[7140] = ~16'b0;
    assign data[7141] = ~16'b0;
    assign data[7142] = ~16'b0;
    assign data[7143] = ~16'b0;
    assign data[7144] = ~16'b0;
    assign data[7145] = ~16'b0;
    assign data[7146] = ~16'b0;
    assign data[7147] = ~16'b0;
    assign data[7148] = ~16'b0;
    assign data[7149] = ~16'b0;
    assign data[7150] = ~16'b0;
    assign data[7151] = ~16'b0;
    assign data[7152] = ~16'b0;
    assign data[7153] = ~16'b0;
    assign data[7154] = ~16'b0;
    assign data[7155] = ~16'b0;
    assign data[7156] = ~16'b0;
    assign data[7157] = ~16'b0;
    assign data[7158] = ~16'b0;
    assign data[7159] = ~16'b0;
    assign data[7160] = ~16'b0;
    assign data[7161] = ~16'b0;
    assign data[7162] = ~16'b0;
    assign data[7163] = ~16'b0;
    assign data[7164] = ~16'b0;
    assign data[7165] = ~16'b0;
    assign data[7166] = ~16'b0;
    assign data[7167] = ~16'b0;
    assign data[7168] = ~16'b0;
    assign data[7169] = ~16'b0;
    assign data[7170] = ~16'b0;
    assign data[7171] = ~16'b0;
    assign data[7172] = ~16'b0;
    assign data[7173] = ~16'b0;
    assign data[7174] = ~16'b0;
    assign data[7175] = ~16'b0;
    assign data[7176] = ~16'b0;
    assign data[7177] = ~16'b0;
    assign data[7178] = ~16'b0;
    assign data[7179] = ~16'b0;
    assign data[7180] = ~16'b0;
    assign data[7181] = ~16'b0;
    assign data[7182] = ~16'b0;
    assign data[7183] = ~16'b0;
    assign data[7184] = ~16'b0;
    assign data[7185] = ~16'b0;
    assign data[7186] = ~16'b0;
    assign data[7187] = ~16'b0;
    assign data[7188] = ~16'b0;
    assign data[7189] = ~16'b0;
    assign data[7190] = ~16'b0;
    assign data[7191] = ~16'b0;
    assign data[7192] = ~16'b0;
    assign data[7193] = ~16'b0;
    assign data[7194] = ~16'b0;
    assign data[7195] = ~16'b0;
    assign data[7196] = ~16'b0;
    assign data[7197] = ~16'b0;
    assign data[7198] = ~16'b0;
    assign data[7199] = ~16'b0;
    assign data[7200] = ~16'b0;
    assign data[7201] = ~16'b0;
    assign data[7202] = ~16'b0;
    assign data[7203] = ~16'b0;
    assign data[7204] = ~16'b0;
    assign data[7205] = ~16'b0;
    assign data[7206] = ~16'b0;
    assign data[7207] = ~16'b0;
    assign data[7208] = ~16'b0;
    assign data[7209] = ~16'b0;
    assign data[7210] = ~16'b0;
    assign data[7211] = ~16'b0;
    assign data[7212] = ~16'b0;
    assign data[7213] = ~16'b0;
    assign data[7214] = ~16'b0;
    assign data[7215] = ~16'b0;
    assign data[7216] = ~16'b0;
    assign data[7217] = ~16'b0;
    assign data[7218] = ~16'b0;
    assign data[7219] = ~16'b0;
    assign data[7220] = ~16'b0;
    assign data[7221] = ~16'b0;
    assign data[7222] = ~16'b0;
    assign data[7223] = ~16'b0;
    assign data[7224] = ~16'b0;
    assign data[7225] = ~16'b0;
    assign data[7226] = ~16'b0;
    assign data[7227] = ~16'b0;
    assign data[7228] = ~16'b0;
    assign data[7229] = ~16'b0;
    assign data[7230] = ~16'b0;
    assign data[7231] = ~16'b0;
    assign data[7232] = ~16'b0;
    assign data[7233] = ~16'b0;
    assign data[7234] = ~16'b0;
    assign data[7235] = ~16'b0;
    assign data[7236] = ~16'b0;
    assign data[7237] = ~16'b0;
    assign data[7238] = ~16'b0;
    assign data[7239] = ~16'b0;
    assign data[7240] = ~16'b0;
    assign data[7241] = ~16'b0;
    assign data[7242] = ~16'b0;
    assign data[7243] = ~16'b0;
    assign data[7244] = ~16'b0;
    assign data[7245] = ~16'b0;
    assign data[7246] = ~16'b0;
    assign data[7247] = ~16'b0;
    assign data[7248] = ~16'b0;
    assign data[7249] = ~16'b0;
    assign data[7250] = ~16'b0;
    assign data[7251] = ~16'b0;
    assign data[7252] = ~16'b0;
    assign data[7253] = ~16'b0;
    assign data[7254] = ~16'b0;
    assign data[7255] = ~16'b0;
    assign data[7256] = ~16'b0;
    assign data[7257] = ~16'b0;
    assign data[7258] = ~16'b0;
    assign data[7259] = ~16'b0;
    assign data[7260] = ~16'b0;
    assign data[7261] = ~16'b0;
    assign data[7262] = ~16'b0;
    assign data[7263] = ~16'b0;
    assign data[7264] = ~16'b0;
    assign data[7265] = ~16'b0;
    assign data[7266] = ~16'b0;
    assign data[7267] = ~16'b0;
    assign data[7268] = ~16'b0;
    assign data[7269] = ~16'b0;
    assign data[7270] = ~16'b0;
    assign data[7271] = ~16'b0;
    assign data[7272] = ~16'b0;
    assign data[7273] = ~16'b0;
    assign data[7274] = ~16'b0;
    assign data[7275] = ~16'b0;
    assign data[7276] = ~16'b0;
    assign data[7277] = ~16'b0;
    assign data[7278] = ~16'b0;
    assign data[7279] = ~16'b0;
    assign data[7280] = ~16'b0;
    assign data[7281] = ~16'b0;
    assign data[7282] = ~16'b0;
    assign data[7283] = ~16'b0;
    assign data[7284] = ~16'b0;
    assign data[7285] = ~16'b0;
    assign data[7286] = ~16'b0;
    assign data[7287] = ~16'b0;
    assign data[7288] = ~16'b0;
    assign data[7289] = ~16'b0;
    assign data[7290] = ~16'b0;
    assign data[7291] = ~16'b0;
    assign data[7292] = ~16'b0;
    assign data[7293] = ~16'b0;
    assign data[7294] = ~16'b0;
    assign data[7295] = ~16'b0;
    assign data[7296] = ~16'b0;
    assign data[7297] = ~16'b0;
    assign data[7298] = ~16'b0;
    assign data[7299] = ~16'b0;
    assign data[7300] = ~16'b0;
    assign data[7301] = ~16'b0;
    assign data[7302] = ~16'b0;
    assign data[7303] = ~16'b0;
    assign data[7304] = ~16'b0;
    assign data[7305] = ~16'b0;
    assign data[7306] = ~16'b0;
    assign data[7307] = ~16'b0;
    assign data[7308] = ~16'b0;
    assign data[7309] = ~16'b0;
    assign data[7310] = ~16'b0;
    assign data[7311] = ~16'b0;
    assign data[7312] = ~16'b0;
    assign data[7313] = ~16'b0;
    assign data[7314] = ~16'b0;
    assign data[7315] = ~16'b0;
    assign data[7316] = ~16'b0;
    assign data[7317] = ~16'b0;
    assign data[7318] = ~16'b0;
    assign data[7319] = ~16'b0;
    assign data[7320] = ~16'b0;
    assign data[7321] = ~16'b0;
    assign data[7322] = ~16'b0;
    assign data[7323] = ~16'b0;
    assign data[7324] = ~16'b0;
    assign data[7325] = ~16'b0;
    assign data[7326] = ~16'b0;
    assign data[7327] = ~16'b0;
    assign data[7328] = ~16'b0;
    assign data[7329] = ~16'b0;
    assign data[7330] = ~16'b0;
    assign data[7331] = ~16'b0;
    assign data[7332] = ~16'b0;
    assign data[7333] = ~16'b0;
    assign data[7334] = ~16'b0;
    assign data[7335] = ~16'b0;
    assign data[7336] = ~16'b0;
    assign data[7337] = ~16'b0;
    assign data[7338] = ~16'b0;
    assign data[7339] = ~16'b0;
    assign data[7340] = ~16'b0;
    assign data[7341] = ~16'b0;
    assign data[7342] = ~16'b0;
    assign data[7343] = ~16'b0;
    assign data[7344] = ~16'b0;
    assign data[7345] = ~16'b0;
    assign data[7346] = ~16'b0;
    assign data[7347] = ~16'b0;
    assign data[7348] = ~16'b0;
    assign data[7349] = ~16'b0;
    assign data[7350] = ~16'b0;
    assign data[7351] = ~16'b0;
    assign data[7352] = ~16'b0;
    assign data[7353] = ~16'b0;
    assign data[7354] = ~16'b0;
    assign data[7355] = ~16'b0;
    assign data[7356] = ~16'b0;
    assign data[7357] = ~16'b0;
    assign data[7358] = ~16'b0;
    assign data[7359] = ~16'b0;
    assign data[7360] = ~16'b0;
    assign data[7361] = ~16'b0;
    assign data[7362] = ~16'b0;
    assign data[7363] = ~16'b0;
    assign data[7364] = ~16'b0;
    assign data[7365] = ~16'b0;
    assign data[7366] = ~16'b0;
    assign data[7367] = ~16'b0;
    assign data[7368] = ~16'b0;
    assign data[7369] = ~16'b0;
    assign data[7370] = ~16'b0;
    assign data[7371] = ~16'b0;
    assign data[7372] = ~16'b0;
    assign data[7373] = ~16'b0;
    assign data[7374] = ~16'b0;
    assign data[7375] = ~16'b0;
    assign data[7376] = ~16'b0;
    assign data[7377] = ~16'b0;
    assign data[7378] = ~16'b0;
    assign data[7379] = ~16'b0;
    

endmodule


